module wallace_tree( 
    input clk,
    input rst_n,
    input [131:0] x_0,
input [131:0] x_1,
input [131:0] x_2,
input [131:0] x_3,
input [131:0] x_4,
input [131:0] x_5,
input [131:0] x_6,
input [131:0] x_7,
input [131:0] x_8,
input [131:0] x_9,
input [131:0] x_10,
input [131:0] x_11,
input [131:0] x_12,
input [131:0] x_13,
input [131:0] x_14,
input [131:0] x_15,
input [131:0] x_16,
input [131:0] x_17,
input [131:0] x_18,
input [131:0] x_19,
input [131:0] x_20,
input [131:0] x_21,
input [131:0] x_22,
input [131:0] x_23,
input [131:0] x_24,
input [131:0] x_25,
input [131:0] x_26,
input [131:0] x_27,
input [131:0] x_28,
input [131:0] x_29,
input [131:0] x_30,
input [131:0] x_31,
input [131:0] x_32,

output [131:0] c,
output [131:0] s,
 input [31:0] c_last_bit_0
);
wire [31:0] c_in_0;
wire [31:0] c_in_1;
wire [31:0] c_in_2;
wire [31:0] c_in_3;
wire [31:0] c_in_4;
wire [31:0] c_in_5;
wire [31:0] c_in_6;
wire [31:0] c_in_7;
wire [31:0] c_in_8;
wire [31:0] c_in_9;
wire [31:0] c_in_10;
wire [31:0] c_in_11;
wire [31:0] c_in_12;
wire [31:0] c_in_13;
wire [31:0] c_in_14;
wire [31:0] c_in_15;
wire [31:0] c_in_16;
wire [31:0] c_in_17;
wire [31:0] c_in_18;
wire [31:0] c_in_19;
wire [31:0] c_in_20;
wire [31:0] c_in_21;
wire [31:0] c_in_22;
wire [31:0] c_in_23;
wire [31:0] c_in_24;
wire [31:0] c_in_25;
wire [31:0] c_in_26;
wire [31:0] c_in_27;
wire [31:0] c_in_28;
wire [31:0] c_in_29;
wire [31:0] c_in_30;
wire [31:0] c_in_31;
wire [31:0] c_in_32;
wire [31:0] c_in_33;
wire [31:0] c_in_34;
wire [31:0] c_in_35;
wire [31:0] c_in_36;
wire [31:0] c_in_37;
wire [31:0] c_in_38;
wire [31:0] c_in_39;
wire [31:0] c_in_40;
wire [31:0] c_in_41;
wire [31:0] c_in_42;
wire [31:0] c_in_43;
wire [31:0] c_in_44;
wire [31:0] c_in_45;
wire [31:0] c_in_46;
wire [31:0] c_in_47;
wire [31:0] c_in_48;
wire [31:0] c_in_49;
wire [31:0] c_in_50;
wire [31:0] c_in_51;
wire [31:0] c_in_52;
wire [31:0] c_in_53;
wire [31:0] c_in_54;
wire [31:0] c_in_55;
wire [31:0] c_in_56;
wire [31:0] c_in_57;
wire [31:0] c_in_58;
wire [31:0] c_in_59;
wire [31:0] c_in_60;
wire [31:0] c_in_61;
wire [31:0] c_in_62;
wire [31:0] c_in_63;
wire [31:0] c_in_64;
wire [31:0] c_in_65;
wire [31:0] c_in_66;
wire [31:0] c_in_67;
wire [31:0] c_in_68;
wire [31:0] c_in_69;
wire [31:0] c_in_70;
wire [31:0] c_in_71;
wire [31:0] c_in_72;
wire [31:0] c_in_73;
wire [31:0] c_in_74;
wire [31:0] c_in_75;
wire [31:0] c_in_76;
wire [31:0] c_in_77;
wire [31:0] c_in_78;
wire [31:0] c_in_79;
wire [31:0] c_in_80;
wire [31:0] c_in_81;
wire [31:0] c_in_82;
wire [31:0] c_in_83;
wire [31:0] c_in_84;
wire [31:0] c_in_85;
wire [31:0] c_in_86;
wire [31:0] c_in_87;
wire [31:0] c_in_88;
wire [31:0] c_in_89;
wire [31:0] c_in_90;
wire [31:0] c_in_91;
wire [31:0] c_in_92;
wire [31:0] c_in_93;
wire [31:0] c_in_94;
wire [31:0] c_in_95;
wire [31:0] c_in_96;
wire [31:0] c_in_97;
wire [31:0] c_in_98;
wire [31:0] c_in_99;
wire [31:0] c_in_100;
wire [31:0] c_in_101;
wire [31:0] c_in_102;
wire [31:0] c_in_103;
wire [31:0] c_in_104;
wire [31:0] c_in_105;
wire [31:0] c_in_106;
wire [31:0] c_in_107;
wire [31:0] c_in_108;
wire [31:0] c_in_109;
wire [31:0] c_in_110;
wire [31:0] c_in_111;
wire [31:0] c_in_112;
wire [31:0] c_in_113;
wire [31:0] c_in_114;
wire [31:0] c_in_115;
wire [31:0] c_in_116;
wire [31:0] c_in_117;
wire [31:0] c_in_118;
wire [31:0] c_in_119;
wire [31:0] c_in_120;
wire [31:0] c_in_121;
wire [31:0] c_in_122;
wire [31:0] c_in_123;
wire [31:0] c_in_124;
wire [31:0] c_in_125;
wire [31:0] c_in_126;
wire [31:0] c_in_127;
wire [31:0] c_in_128;
wire [31:0] c_in_129;
wire [31:0] c_in_130;
wire [31:0] c_in_131;
assign c_in_0 = c_last_bit_0;
wire  c_0;
wire  s_0;
wallace_tree_ w0(.clk(clk),.rst_n(rst_n),.a({x_0[0],x_1[0],x_2[0],x_3[0],x_4[0],x_5[0],x_6[0],x_7[0],x_8[0],x_9[0],x_10[0],x_11[0],x_12[0],x_13[0],x_14[0],x_15[0],x_16[0],x_17[0],x_18[0],x_19[0],x_20[0],x_21[0],x_22[0],x_23[0],x_24[0],x_25[0],x_26[0],x_27[0],x_28[0],x_29[0],x_30[0],x_31[0],x_32[0]}),.c_in(c_in_0),.c_out(c_in_1),.s(s_0),.c(c_0));
wire  c_1;
wire  s_1;
wallace_tree_ w1(.clk(clk),.rst_n(rst_n),.a({x_0[1],x_1[1],x_2[1],x_3[1],x_4[1],x_5[1],x_6[1],x_7[1],x_8[1],x_9[1],x_10[1],x_11[1],x_12[1],x_13[1],x_14[1],x_15[1],x_16[1],x_17[1],x_18[1],x_19[1],x_20[1],x_21[1],x_22[1],x_23[1],x_24[1],x_25[1],x_26[1],x_27[1],x_28[1],x_29[1],x_30[1],x_31[1],x_32[1]}),.c_in(c_in_1),.c_out(c_in_2),.s(s_1),.c(c_1));
wire  c_2;
wire  s_2;
wallace_tree_ w2(.clk(clk),.rst_n(rst_n),.a({x_0[2],x_1[2],x_2[2],x_3[2],x_4[2],x_5[2],x_6[2],x_7[2],x_8[2],x_9[2],x_10[2],x_11[2],x_12[2],x_13[2],x_14[2],x_15[2],x_16[2],x_17[2],x_18[2],x_19[2],x_20[2],x_21[2],x_22[2],x_23[2],x_24[2],x_25[2],x_26[2],x_27[2],x_28[2],x_29[2],x_30[2],x_31[2],x_32[2]}),.c_in(c_in_2),.c_out(c_in_3),.s(s_2),.c(c_2));
wire  c_3;
wire  s_3;
wallace_tree_ w3(.clk(clk),.rst_n(rst_n),.a({x_0[3],x_1[3],x_2[3],x_3[3],x_4[3],x_5[3],x_6[3],x_7[3],x_8[3],x_9[3],x_10[3],x_11[3],x_12[3],x_13[3],x_14[3],x_15[3],x_16[3],x_17[3],x_18[3],x_19[3],x_20[3],x_21[3],x_22[3],x_23[3],x_24[3],x_25[3],x_26[3],x_27[3],x_28[3],x_29[3],x_30[3],x_31[3],x_32[3]}),.c_in(c_in_3),.c_out(c_in_4),.s(s_3),.c(c_3));
wire  c_4;
wire  s_4;
wallace_tree_ w4(.clk(clk),.rst_n(rst_n),.a({x_0[4],x_1[4],x_2[4],x_3[4],x_4[4],x_5[4],x_6[4],x_7[4],x_8[4],x_9[4],x_10[4],x_11[4],x_12[4],x_13[4],x_14[4],x_15[4],x_16[4],x_17[4],x_18[4],x_19[4],x_20[4],x_21[4],x_22[4],x_23[4],x_24[4],x_25[4],x_26[4],x_27[4],x_28[4],x_29[4],x_30[4],x_31[4],x_32[4]}),.c_in(c_in_4),.c_out(c_in_5),.s(s_4),.c(c_4));
wire  c_5;
wire  s_5;
wallace_tree_ w5(.clk(clk),.rst_n(rst_n),.a({x_0[5],x_1[5],x_2[5],x_3[5],x_4[5],x_5[5],x_6[5],x_7[5],x_8[5],x_9[5],x_10[5],x_11[5],x_12[5],x_13[5],x_14[5],x_15[5],x_16[5],x_17[5],x_18[5],x_19[5],x_20[5],x_21[5],x_22[5],x_23[5],x_24[5],x_25[5],x_26[5],x_27[5],x_28[5],x_29[5],x_30[5],x_31[5],x_32[5]}),.c_in(c_in_5),.c_out(c_in_6),.s(s_5),.c(c_5));
wire  c_6;
wire  s_6;
wallace_tree_ w6(.clk(clk),.rst_n(rst_n),.a({x_0[6],x_1[6],x_2[6],x_3[6],x_4[6],x_5[6],x_6[6],x_7[6],x_8[6],x_9[6],x_10[6],x_11[6],x_12[6],x_13[6],x_14[6],x_15[6],x_16[6],x_17[6],x_18[6],x_19[6],x_20[6],x_21[6],x_22[6],x_23[6],x_24[6],x_25[6],x_26[6],x_27[6],x_28[6],x_29[6],x_30[6],x_31[6],x_32[6]}),.c_in(c_in_6),.c_out(c_in_7),.s(s_6),.c(c_6));
wire  c_7;
wire  s_7;
wallace_tree_ w7(.clk(clk),.rst_n(rst_n),.a({x_0[7],x_1[7],x_2[7],x_3[7],x_4[7],x_5[7],x_6[7],x_7[7],x_8[7],x_9[7],x_10[7],x_11[7],x_12[7],x_13[7],x_14[7],x_15[7],x_16[7],x_17[7],x_18[7],x_19[7],x_20[7],x_21[7],x_22[7],x_23[7],x_24[7],x_25[7],x_26[7],x_27[7],x_28[7],x_29[7],x_30[7],x_31[7],x_32[7]}),.c_in(c_in_7),.c_out(c_in_8),.s(s_7),.c(c_7));
wire  c_8;
wire  s_8;
wallace_tree_ w8(.clk(clk),.rst_n(rst_n),.a({x_0[8],x_1[8],x_2[8],x_3[8],x_4[8],x_5[8],x_6[8],x_7[8],x_8[8],x_9[8],x_10[8],x_11[8],x_12[8],x_13[8],x_14[8],x_15[8],x_16[8],x_17[8],x_18[8],x_19[8],x_20[8],x_21[8],x_22[8],x_23[8],x_24[8],x_25[8],x_26[8],x_27[8],x_28[8],x_29[8],x_30[8],x_31[8],x_32[8]}),.c_in(c_in_8),.c_out(c_in_9),.s(s_8),.c(c_8));
wire  c_9;
wire  s_9;
wallace_tree_ w9(.clk(clk),.rst_n(rst_n),.a({x_0[9],x_1[9],x_2[9],x_3[9],x_4[9],x_5[9],x_6[9],x_7[9],x_8[9],x_9[9],x_10[9],x_11[9],x_12[9],x_13[9],x_14[9],x_15[9],x_16[9],x_17[9],x_18[9],x_19[9],x_20[9],x_21[9],x_22[9],x_23[9],x_24[9],x_25[9],x_26[9],x_27[9],x_28[9],x_29[9],x_30[9],x_31[9],x_32[9]}),.c_in(c_in_9),.c_out(c_in_10),.s(s_9),.c(c_9));
wire  c_10;
wire  s_10;
wallace_tree_ w10(.clk(clk),.rst_n(rst_n),.a({x_0[10],x_1[10],x_2[10],x_3[10],x_4[10],x_5[10],x_6[10],x_7[10],x_8[10],x_9[10],x_10[10],x_11[10],x_12[10],x_13[10],x_14[10],x_15[10],x_16[10],x_17[10],x_18[10],x_19[10],x_20[10],x_21[10],x_22[10],x_23[10],x_24[10],x_25[10],x_26[10],x_27[10],x_28[10],x_29[10],x_30[10],x_31[10],x_32[10]}),.c_in(c_in_10),.c_out(c_in_11),.s(s_10),.c(c_10));
wire  c_11;
wire  s_11;
wallace_tree_ w11(.clk(clk),.rst_n(rst_n),.a({x_0[11],x_1[11],x_2[11],x_3[11],x_4[11],x_5[11],x_6[11],x_7[11],x_8[11],x_9[11],x_10[11],x_11[11],x_12[11],x_13[11],x_14[11],x_15[11],x_16[11],x_17[11],x_18[11],x_19[11],x_20[11],x_21[11],x_22[11],x_23[11],x_24[11],x_25[11],x_26[11],x_27[11],x_28[11],x_29[11],x_30[11],x_31[11],x_32[11]}),.c_in(c_in_11),.c_out(c_in_12),.s(s_11),.c(c_11));
wire  c_12;
wire  s_12;
wallace_tree_ w12(.clk(clk),.rst_n(rst_n),.a({x_0[12],x_1[12],x_2[12],x_3[12],x_4[12],x_5[12],x_6[12],x_7[12],x_8[12],x_9[12],x_10[12],x_11[12],x_12[12],x_13[12],x_14[12],x_15[12],x_16[12],x_17[12],x_18[12],x_19[12],x_20[12],x_21[12],x_22[12],x_23[12],x_24[12],x_25[12],x_26[12],x_27[12],x_28[12],x_29[12],x_30[12],x_31[12],x_32[12]}),.c_in(c_in_12),.c_out(c_in_13),.s(s_12),.c(c_12));
wire  c_13;
wire  s_13;
wallace_tree_ w13(.clk(clk),.rst_n(rst_n),.a({x_0[13],x_1[13],x_2[13],x_3[13],x_4[13],x_5[13],x_6[13],x_7[13],x_8[13],x_9[13],x_10[13],x_11[13],x_12[13],x_13[13],x_14[13],x_15[13],x_16[13],x_17[13],x_18[13],x_19[13],x_20[13],x_21[13],x_22[13],x_23[13],x_24[13],x_25[13],x_26[13],x_27[13],x_28[13],x_29[13],x_30[13],x_31[13],x_32[13]}),.c_in(c_in_13),.c_out(c_in_14),.s(s_13),.c(c_13));
wire  c_14;
wire  s_14;
wallace_tree_ w14(.clk(clk),.rst_n(rst_n),.a({x_0[14],x_1[14],x_2[14],x_3[14],x_4[14],x_5[14],x_6[14],x_7[14],x_8[14],x_9[14],x_10[14],x_11[14],x_12[14],x_13[14],x_14[14],x_15[14],x_16[14],x_17[14],x_18[14],x_19[14],x_20[14],x_21[14],x_22[14],x_23[14],x_24[14],x_25[14],x_26[14],x_27[14],x_28[14],x_29[14],x_30[14],x_31[14],x_32[14]}),.c_in(c_in_14),.c_out(c_in_15),.s(s_14),.c(c_14));
wire  c_15;
wire  s_15;
wallace_tree_ w15(.clk(clk),.rst_n(rst_n),.a({x_0[15],x_1[15],x_2[15],x_3[15],x_4[15],x_5[15],x_6[15],x_7[15],x_8[15],x_9[15],x_10[15],x_11[15],x_12[15],x_13[15],x_14[15],x_15[15],x_16[15],x_17[15],x_18[15],x_19[15],x_20[15],x_21[15],x_22[15],x_23[15],x_24[15],x_25[15],x_26[15],x_27[15],x_28[15],x_29[15],x_30[15],x_31[15],x_32[15]}),.c_in(c_in_15),.c_out(c_in_16),.s(s_15),.c(c_15));
wire  c_16;
wire  s_16;
wallace_tree_ w16(.clk(clk),.rst_n(rst_n),.a({x_0[16],x_1[16],x_2[16],x_3[16],x_4[16],x_5[16],x_6[16],x_7[16],x_8[16],x_9[16],x_10[16],x_11[16],x_12[16],x_13[16],x_14[16],x_15[16],x_16[16],x_17[16],x_18[16],x_19[16],x_20[16],x_21[16],x_22[16],x_23[16],x_24[16],x_25[16],x_26[16],x_27[16],x_28[16],x_29[16],x_30[16],x_31[16],x_32[16]}),.c_in(c_in_16),.c_out(c_in_17),.s(s_16),.c(c_16));
wire  c_17;
wire  s_17;
wallace_tree_ w17(.clk(clk),.rst_n(rst_n),.a({x_0[17],x_1[17],x_2[17],x_3[17],x_4[17],x_5[17],x_6[17],x_7[17],x_8[17],x_9[17],x_10[17],x_11[17],x_12[17],x_13[17],x_14[17],x_15[17],x_16[17],x_17[17],x_18[17],x_19[17],x_20[17],x_21[17],x_22[17],x_23[17],x_24[17],x_25[17],x_26[17],x_27[17],x_28[17],x_29[17],x_30[17],x_31[17],x_32[17]}),.c_in(c_in_17),.c_out(c_in_18),.s(s_17),.c(c_17));
wire  c_18;
wire  s_18;
wallace_tree_ w18(.clk(clk),.rst_n(rst_n),.a({x_0[18],x_1[18],x_2[18],x_3[18],x_4[18],x_5[18],x_6[18],x_7[18],x_8[18],x_9[18],x_10[18],x_11[18],x_12[18],x_13[18],x_14[18],x_15[18],x_16[18],x_17[18],x_18[18],x_19[18],x_20[18],x_21[18],x_22[18],x_23[18],x_24[18],x_25[18],x_26[18],x_27[18],x_28[18],x_29[18],x_30[18],x_31[18],x_32[18]}),.c_in(c_in_18),.c_out(c_in_19),.s(s_18),.c(c_18));
wire  c_19;
wire  s_19;
wallace_tree_ w19(.clk(clk),.rst_n(rst_n),.a({x_0[19],x_1[19],x_2[19],x_3[19],x_4[19],x_5[19],x_6[19],x_7[19],x_8[19],x_9[19],x_10[19],x_11[19],x_12[19],x_13[19],x_14[19],x_15[19],x_16[19],x_17[19],x_18[19],x_19[19],x_20[19],x_21[19],x_22[19],x_23[19],x_24[19],x_25[19],x_26[19],x_27[19],x_28[19],x_29[19],x_30[19],x_31[19],x_32[19]}),.c_in(c_in_19),.c_out(c_in_20),.s(s_19),.c(c_19));
wire  c_20;
wire  s_20;
wallace_tree_ w20(.clk(clk),.rst_n(rst_n),.a({x_0[20],x_1[20],x_2[20],x_3[20],x_4[20],x_5[20],x_6[20],x_7[20],x_8[20],x_9[20],x_10[20],x_11[20],x_12[20],x_13[20],x_14[20],x_15[20],x_16[20],x_17[20],x_18[20],x_19[20],x_20[20],x_21[20],x_22[20],x_23[20],x_24[20],x_25[20],x_26[20],x_27[20],x_28[20],x_29[20],x_30[20],x_31[20],x_32[20]}),.c_in(c_in_20),.c_out(c_in_21),.s(s_20),.c(c_20));
wire  c_21;
wire  s_21;
wallace_tree_ w21(.clk(clk),.rst_n(rst_n),.a({x_0[21],x_1[21],x_2[21],x_3[21],x_4[21],x_5[21],x_6[21],x_7[21],x_8[21],x_9[21],x_10[21],x_11[21],x_12[21],x_13[21],x_14[21],x_15[21],x_16[21],x_17[21],x_18[21],x_19[21],x_20[21],x_21[21],x_22[21],x_23[21],x_24[21],x_25[21],x_26[21],x_27[21],x_28[21],x_29[21],x_30[21],x_31[21],x_32[21]}),.c_in(c_in_21),.c_out(c_in_22),.s(s_21),.c(c_21));
wire  c_22;
wire  s_22;
wallace_tree_ w22(.clk(clk),.rst_n(rst_n),.a({x_0[22],x_1[22],x_2[22],x_3[22],x_4[22],x_5[22],x_6[22],x_7[22],x_8[22],x_9[22],x_10[22],x_11[22],x_12[22],x_13[22],x_14[22],x_15[22],x_16[22],x_17[22],x_18[22],x_19[22],x_20[22],x_21[22],x_22[22],x_23[22],x_24[22],x_25[22],x_26[22],x_27[22],x_28[22],x_29[22],x_30[22],x_31[22],x_32[22]}),.c_in(c_in_22),.c_out(c_in_23),.s(s_22),.c(c_22));
wire  c_23;
wire  s_23;
wallace_tree_ w23(.clk(clk),.rst_n(rst_n),.a({x_0[23],x_1[23],x_2[23],x_3[23],x_4[23],x_5[23],x_6[23],x_7[23],x_8[23],x_9[23],x_10[23],x_11[23],x_12[23],x_13[23],x_14[23],x_15[23],x_16[23],x_17[23],x_18[23],x_19[23],x_20[23],x_21[23],x_22[23],x_23[23],x_24[23],x_25[23],x_26[23],x_27[23],x_28[23],x_29[23],x_30[23],x_31[23],x_32[23]}),.c_in(c_in_23),.c_out(c_in_24),.s(s_23),.c(c_23));
wire  c_24;
wire  s_24;
wallace_tree_ w24(.clk(clk),.rst_n(rst_n),.a({x_0[24],x_1[24],x_2[24],x_3[24],x_4[24],x_5[24],x_6[24],x_7[24],x_8[24],x_9[24],x_10[24],x_11[24],x_12[24],x_13[24],x_14[24],x_15[24],x_16[24],x_17[24],x_18[24],x_19[24],x_20[24],x_21[24],x_22[24],x_23[24],x_24[24],x_25[24],x_26[24],x_27[24],x_28[24],x_29[24],x_30[24],x_31[24],x_32[24]}),.c_in(c_in_24),.c_out(c_in_25),.s(s_24),.c(c_24));
wire  c_25;
wire  s_25;
wallace_tree_ w25(.clk(clk),.rst_n(rst_n),.a({x_0[25],x_1[25],x_2[25],x_3[25],x_4[25],x_5[25],x_6[25],x_7[25],x_8[25],x_9[25],x_10[25],x_11[25],x_12[25],x_13[25],x_14[25],x_15[25],x_16[25],x_17[25],x_18[25],x_19[25],x_20[25],x_21[25],x_22[25],x_23[25],x_24[25],x_25[25],x_26[25],x_27[25],x_28[25],x_29[25],x_30[25],x_31[25],x_32[25]}),.c_in(c_in_25),.c_out(c_in_26),.s(s_25),.c(c_25));
wire  c_26;
wire  s_26;
wallace_tree_ w26(.clk(clk),.rst_n(rst_n),.a({x_0[26],x_1[26],x_2[26],x_3[26],x_4[26],x_5[26],x_6[26],x_7[26],x_8[26],x_9[26],x_10[26],x_11[26],x_12[26],x_13[26],x_14[26],x_15[26],x_16[26],x_17[26],x_18[26],x_19[26],x_20[26],x_21[26],x_22[26],x_23[26],x_24[26],x_25[26],x_26[26],x_27[26],x_28[26],x_29[26],x_30[26],x_31[26],x_32[26]}),.c_in(c_in_26),.c_out(c_in_27),.s(s_26),.c(c_26));
wire  c_27;
wire  s_27;
wallace_tree_ w27(.clk(clk),.rst_n(rst_n),.a({x_0[27],x_1[27],x_2[27],x_3[27],x_4[27],x_5[27],x_6[27],x_7[27],x_8[27],x_9[27],x_10[27],x_11[27],x_12[27],x_13[27],x_14[27],x_15[27],x_16[27],x_17[27],x_18[27],x_19[27],x_20[27],x_21[27],x_22[27],x_23[27],x_24[27],x_25[27],x_26[27],x_27[27],x_28[27],x_29[27],x_30[27],x_31[27],x_32[27]}),.c_in(c_in_27),.c_out(c_in_28),.s(s_27),.c(c_27));
wire  c_28;
wire  s_28;
wallace_tree_ w28(.clk(clk),.rst_n(rst_n),.a({x_0[28],x_1[28],x_2[28],x_3[28],x_4[28],x_5[28],x_6[28],x_7[28],x_8[28],x_9[28],x_10[28],x_11[28],x_12[28],x_13[28],x_14[28],x_15[28],x_16[28],x_17[28],x_18[28],x_19[28],x_20[28],x_21[28],x_22[28],x_23[28],x_24[28],x_25[28],x_26[28],x_27[28],x_28[28],x_29[28],x_30[28],x_31[28],x_32[28]}),.c_in(c_in_28),.c_out(c_in_29),.s(s_28),.c(c_28));
wire  c_29;
wire  s_29;
wallace_tree_ w29(.clk(clk),.rst_n(rst_n),.a({x_0[29],x_1[29],x_2[29],x_3[29],x_4[29],x_5[29],x_6[29],x_7[29],x_8[29],x_9[29],x_10[29],x_11[29],x_12[29],x_13[29],x_14[29],x_15[29],x_16[29],x_17[29],x_18[29],x_19[29],x_20[29],x_21[29],x_22[29],x_23[29],x_24[29],x_25[29],x_26[29],x_27[29],x_28[29],x_29[29],x_30[29],x_31[29],x_32[29]}),.c_in(c_in_29),.c_out(c_in_30),.s(s_29),.c(c_29));
wire  c_30;
wire  s_30;
wallace_tree_ w30(.clk(clk),.rst_n(rst_n),.a({x_0[30],x_1[30],x_2[30],x_3[30],x_4[30],x_5[30],x_6[30],x_7[30],x_8[30],x_9[30],x_10[30],x_11[30],x_12[30],x_13[30],x_14[30],x_15[30],x_16[30],x_17[30],x_18[30],x_19[30],x_20[30],x_21[30],x_22[30],x_23[30],x_24[30],x_25[30],x_26[30],x_27[30],x_28[30],x_29[30],x_30[30],x_31[30],x_32[30]}),.c_in(c_in_30),.c_out(c_in_31),.s(s_30),.c(c_30));
wire  c_31;
wire  s_31;
wallace_tree_ w31(.clk(clk),.rst_n(rst_n),.a({x_0[31],x_1[31],x_2[31],x_3[31],x_4[31],x_5[31],x_6[31],x_7[31],x_8[31],x_9[31],x_10[31],x_11[31],x_12[31],x_13[31],x_14[31],x_15[31],x_16[31],x_17[31],x_18[31],x_19[31],x_20[31],x_21[31],x_22[31],x_23[31],x_24[31],x_25[31],x_26[31],x_27[31],x_28[31],x_29[31],x_30[31],x_31[31],x_32[31]}),.c_in(c_in_31),.c_out(c_in_32),.s(s_31),.c(c_31));
wire  c_32;
wire  s_32;
wallace_tree_ w32(.clk(clk),.rst_n(rst_n),.a({x_0[32],x_1[32],x_2[32],x_3[32],x_4[32],x_5[32],x_6[32],x_7[32],x_8[32],x_9[32],x_10[32],x_11[32],x_12[32],x_13[32],x_14[32],x_15[32],x_16[32],x_17[32],x_18[32],x_19[32],x_20[32],x_21[32],x_22[32],x_23[32],x_24[32],x_25[32],x_26[32],x_27[32],x_28[32],x_29[32],x_30[32],x_31[32],x_32[32]}),.c_in(c_in_32),.c_out(c_in_33),.s(s_32),.c(c_32));
wire  c_33;
wire  s_33;
wallace_tree_ w33(.clk(clk),.rst_n(rst_n),.a({x_0[33],x_1[33],x_2[33],x_3[33],x_4[33],x_5[33],x_6[33],x_7[33],x_8[33],x_9[33],x_10[33],x_11[33],x_12[33],x_13[33],x_14[33],x_15[33],x_16[33],x_17[33],x_18[33],x_19[33],x_20[33],x_21[33],x_22[33],x_23[33],x_24[33],x_25[33],x_26[33],x_27[33],x_28[33],x_29[33],x_30[33],x_31[33],x_32[33]}),.c_in(c_in_33),.c_out(c_in_34),.s(s_33),.c(c_33));
wire  c_34;
wire  s_34;
wallace_tree_ w34(.clk(clk),.rst_n(rst_n),.a({x_0[34],x_1[34],x_2[34],x_3[34],x_4[34],x_5[34],x_6[34],x_7[34],x_8[34],x_9[34],x_10[34],x_11[34],x_12[34],x_13[34],x_14[34],x_15[34],x_16[34],x_17[34],x_18[34],x_19[34],x_20[34],x_21[34],x_22[34],x_23[34],x_24[34],x_25[34],x_26[34],x_27[34],x_28[34],x_29[34],x_30[34],x_31[34],x_32[34]}),.c_in(c_in_34),.c_out(c_in_35),.s(s_34),.c(c_34));
wire  c_35;
wire  s_35;
wallace_tree_ w35(.clk(clk),.rst_n(rst_n),.a({x_0[35],x_1[35],x_2[35],x_3[35],x_4[35],x_5[35],x_6[35],x_7[35],x_8[35],x_9[35],x_10[35],x_11[35],x_12[35],x_13[35],x_14[35],x_15[35],x_16[35],x_17[35],x_18[35],x_19[35],x_20[35],x_21[35],x_22[35],x_23[35],x_24[35],x_25[35],x_26[35],x_27[35],x_28[35],x_29[35],x_30[35],x_31[35],x_32[35]}),.c_in(c_in_35),.c_out(c_in_36),.s(s_35),.c(c_35));
wire  c_36;
wire  s_36;
wallace_tree_ w36(.clk(clk),.rst_n(rst_n),.a({x_0[36],x_1[36],x_2[36],x_3[36],x_4[36],x_5[36],x_6[36],x_7[36],x_8[36],x_9[36],x_10[36],x_11[36],x_12[36],x_13[36],x_14[36],x_15[36],x_16[36],x_17[36],x_18[36],x_19[36],x_20[36],x_21[36],x_22[36],x_23[36],x_24[36],x_25[36],x_26[36],x_27[36],x_28[36],x_29[36],x_30[36],x_31[36],x_32[36]}),.c_in(c_in_36),.c_out(c_in_37),.s(s_36),.c(c_36));
wire  c_37;
wire  s_37;
wallace_tree_ w37(.clk(clk),.rst_n(rst_n),.a({x_0[37],x_1[37],x_2[37],x_3[37],x_4[37],x_5[37],x_6[37],x_7[37],x_8[37],x_9[37],x_10[37],x_11[37],x_12[37],x_13[37],x_14[37],x_15[37],x_16[37],x_17[37],x_18[37],x_19[37],x_20[37],x_21[37],x_22[37],x_23[37],x_24[37],x_25[37],x_26[37],x_27[37],x_28[37],x_29[37],x_30[37],x_31[37],x_32[37]}),.c_in(c_in_37),.c_out(c_in_38),.s(s_37),.c(c_37));
wire  c_38;
wire  s_38;
wallace_tree_ w38(.clk(clk),.rst_n(rst_n),.a({x_0[38],x_1[38],x_2[38],x_3[38],x_4[38],x_5[38],x_6[38],x_7[38],x_8[38],x_9[38],x_10[38],x_11[38],x_12[38],x_13[38],x_14[38],x_15[38],x_16[38],x_17[38],x_18[38],x_19[38],x_20[38],x_21[38],x_22[38],x_23[38],x_24[38],x_25[38],x_26[38],x_27[38],x_28[38],x_29[38],x_30[38],x_31[38],x_32[38]}),.c_in(c_in_38),.c_out(c_in_39),.s(s_38),.c(c_38));
wire  c_39;
wire  s_39;
wallace_tree_ w39(.clk(clk),.rst_n(rst_n),.a({x_0[39],x_1[39],x_2[39],x_3[39],x_4[39],x_5[39],x_6[39],x_7[39],x_8[39],x_9[39],x_10[39],x_11[39],x_12[39],x_13[39],x_14[39],x_15[39],x_16[39],x_17[39],x_18[39],x_19[39],x_20[39],x_21[39],x_22[39],x_23[39],x_24[39],x_25[39],x_26[39],x_27[39],x_28[39],x_29[39],x_30[39],x_31[39],x_32[39]}),.c_in(c_in_39),.c_out(c_in_40),.s(s_39),.c(c_39));
wire  c_40;
wire  s_40;
wallace_tree_ w40(.clk(clk),.rst_n(rst_n),.a({x_0[40],x_1[40],x_2[40],x_3[40],x_4[40],x_5[40],x_6[40],x_7[40],x_8[40],x_9[40],x_10[40],x_11[40],x_12[40],x_13[40],x_14[40],x_15[40],x_16[40],x_17[40],x_18[40],x_19[40],x_20[40],x_21[40],x_22[40],x_23[40],x_24[40],x_25[40],x_26[40],x_27[40],x_28[40],x_29[40],x_30[40],x_31[40],x_32[40]}),.c_in(c_in_40),.c_out(c_in_41),.s(s_40),.c(c_40));
wire  c_41;
wire  s_41;
wallace_tree_ w41(.clk(clk),.rst_n(rst_n),.a({x_0[41],x_1[41],x_2[41],x_3[41],x_4[41],x_5[41],x_6[41],x_7[41],x_8[41],x_9[41],x_10[41],x_11[41],x_12[41],x_13[41],x_14[41],x_15[41],x_16[41],x_17[41],x_18[41],x_19[41],x_20[41],x_21[41],x_22[41],x_23[41],x_24[41],x_25[41],x_26[41],x_27[41],x_28[41],x_29[41],x_30[41],x_31[41],x_32[41]}),.c_in(c_in_41),.c_out(c_in_42),.s(s_41),.c(c_41));
wire  c_42;
wire  s_42;
wallace_tree_ w42(.clk(clk),.rst_n(rst_n),.a({x_0[42],x_1[42],x_2[42],x_3[42],x_4[42],x_5[42],x_6[42],x_7[42],x_8[42],x_9[42],x_10[42],x_11[42],x_12[42],x_13[42],x_14[42],x_15[42],x_16[42],x_17[42],x_18[42],x_19[42],x_20[42],x_21[42],x_22[42],x_23[42],x_24[42],x_25[42],x_26[42],x_27[42],x_28[42],x_29[42],x_30[42],x_31[42],x_32[42]}),.c_in(c_in_42),.c_out(c_in_43),.s(s_42),.c(c_42));
wire  c_43;
wire  s_43;
wallace_tree_ w43(.clk(clk),.rst_n(rst_n),.a({x_0[43],x_1[43],x_2[43],x_3[43],x_4[43],x_5[43],x_6[43],x_7[43],x_8[43],x_9[43],x_10[43],x_11[43],x_12[43],x_13[43],x_14[43],x_15[43],x_16[43],x_17[43],x_18[43],x_19[43],x_20[43],x_21[43],x_22[43],x_23[43],x_24[43],x_25[43],x_26[43],x_27[43],x_28[43],x_29[43],x_30[43],x_31[43],x_32[43]}),.c_in(c_in_43),.c_out(c_in_44),.s(s_43),.c(c_43));
wire  c_44;
wire  s_44;
wallace_tree_ w44(.clk(clk),.rst_n(rst_n),.a({x_0[44],x_1[44],x_2[44],x_3[44],x_4[44],x_5[44],x_6[44],x_7[44],x_8[44],x_9[44],x_10[44],x_11[44],x_12[44],x_13[44],x_14[44],x_15[44],x_16[44],x_17[44],x_18[44],x_19[44],x_20[44],x_21[44],x_22[44],x_23[44],x_24[44],x_25[44],x_26[44],x_27[44],x_28[44],x_29[44],x_30[44],x_31[44],x_32[44]}),.c_in(c_in_44),.c_out(c_in_45),.s(s_44),.c(c_44));
wire  c_45;
wire  s_45;
wallace_tree_ w45(.clk(clk),.rst_n(rst_n),.a({x_0[45],x_1[45],x_2[45],x_3[45],x_4[45],x_5[45],x_6[45],x_7[45],x_8[45],x_9[45],x_10[45],x_11[45],x_12[45],x_13[45],x_14[45],x_15[45],x_16[45],x_17[45],x_18[45],x_19[45],x_20[45],x_21[45],x_22[45],x_23[45],x_24[45],x_25[45],x_26[45],x_27[45],x_28[45],x_29[45],x_30[45],x_31[45],x_32[45]}),.c_in(c_in_45),.c_out(c_in_46),.s(s_45),.c(c_45));
wire  c_46;
wire  s_46;
wallace_tree_ w46(.clk(clk),.rst_n(rst_n),.a({x_0[46],x_1[46],x_2[46],x_3[46],x_4[46],x_5[46],x_6[46],x_7[46],x_8[46],x_9[46],x_10[46],x_11[46],x_12[46],x_13[46],x_14[46],x_15[46],x_16[46],x_17[46],x_18[46],x_19[46],x_20[46],x_21[46],x_22[46],x_23[46],x_24[46],x_25[46],x_26[46],x_27[46],x_28[46],x_29[46],x_30[46],x_31[46],x_32[46]}),.c_in(c_in_46),.c_out(c_in_47),.s(s_46),.c(c_46));
wire  c_47;
wire  s_47;
wallace_tree_ w47(.clk(clk),.rst_n(rst_n),.a({x_0[47],x_1[47],x_2[47],x_3[47],x_4[47],x_5[47],x_6[47],x_7[47],x_8[47],x_9[47],x_10[47],x_11[47],x_12[47],x_13[47],x_14[47],x_15[47],x_16[47],x_17[47],x_18[47],x_19[47],x_20[47],x_21[47],x_22[47],x_23[47],x_24[47],x_25[47],x_26[47],x_27[47],x_28[47],x_29[47],x_30[47],x_31[47],x_32[47]}),.c_in(c_in_47),.c_out(c_in_48),.s(s_47),.c(c_47));
wire  c_48;
wire  s_48;
wallace_tree_ w48(.clk(clk),.rst_n(rst_n),.a({x_0[48],x_1[48],x_2[48],x_3[48],x_4[48],x_5[48],x_6[48],x_7[48],x_8[48],x_9[48],x_10[48],x_11[48],x_12[48],x_13[48],x_14[48],x_15[48],x_16[48],x_17[48],x_18[48],x_19[48],x_20[48],x_21[48],x_22[48],x_23[48],x_24[48],x_25[48],x_26[48],x_27[48],x_28[48],x_29[48],x_30[48],x_31[48],x_32[48]}),.c_in(c_in_48),.c_out(c_in_49),.s(s_48),.c(c_48));
wire  c_49;
wire  s_49;
wallace_tree_ w49(.clk(clk),.rst_n(rst_n),.a({x_0[49],x_1[49],x_2[49],x_3[49],x_4[49],x_5[49],x_6[49],x_7[49],x_8[49],x_9[49],x_10[49],x_11[49],x_12[49],x_13[49],x_14[49],x_15[49],x_16[49],x_17[49],x_18[49],x_19[49],x_20[49],x_21[49],x_22[49],x_23[49],x_24[49],x_25[49],x_26[49],x_27[49],x_28[49],x_29[49],x_30[49],x_31[49],x_32[49]}),.c_in(c_in_49),.c_out(c_in_50),.s(s_49),.c(c_49));
wire  c_50;
wire  s_50;
wallace_tree_ w50(.clk(clk),.rst_n(rst_n),.a({x_0[50],x_1[50],x_2[50],x_3[50],x_4[50],x_5[50],x_6[50],x_7[50],x_8[50],x_9[50],x_10[50],x_11[50],x_12[50],x_13[50],x_14[50],x_15[50],x_16[50],x_17[50],x_18[50],x_19[50],x_20[50],x_21[50],x_22[50],x_23[50],x_24[50],x_25[50],x_26[50],x_27[50],x_28[50],x_29[50],x_30[50],x_31[50],x_32[50]}),.c_in(c_in_50),.c_out(c_in_51),.s(s_50),.c(c_50));
wire  c_51;
wire  s_51;
wallace_tree_ w51(.clk(clk),.rst_n(rst_n),.a({x_0[51],x_1[51],x_2[51],x_3[51],x_4[51],x_5[51],x_6[51],x_7[51],x_8[51],x_9[51],x_10[51],x_11[51],x_12[51],x_13[51],x_14[51],x_15[51],x_16[51],x_17[51],x_18[51],x_19[51],x_20[51],x_21[51],x_22[51],x_23[51],x_24[51],x_25[51],x_26[51],x_27[51],x_28[51],x_29[51],x_30[51],x_31[51],x_32[51]}),.c_in(c_in_51),.c_out(c_in_52),.s(s_51),.c(c_51));
wire  c_52;
wire  s_52;
wallace_tree_ w52(.clk(clk),.rst_n(rst_n),.a({x_0[52],x_1[52],x_2[52],x_3[52],x_4[52],x_5[52],x_6[52],x_7[52],x_8[52],x_9[52],x_10[52],x_11[52],x_12[52],x_13[52],x_14[52],x_15[52],x_16[52],x_17[52],x_18[52],x_19[52],x_20[52],x_21[52],x_22[52],x_23[52],x_24[52],x_25[52],x_26[52],x_27[52],x_28[52],x_29[52],x_30[52],x_31[52],x_32[52]}),.c_in(c_in_52),.c_out(c_in_53),.s(s_52),.c(c_52));
wire  c_53;
wire  s_53;
wallace_tree_ w53(.clk(clk),.rst_n(rst_n),.a({x_0[53],x_1[53],x_2[53],x_3[53],x_4[53],x_5[53],x_6[53],x_7[53],x_8[53],x_9[53],x_10[53],x_11[53],x_12[53],x_13[53],x_14[53],x_15[53],x_16[53],x_17[53],x_18[53],x_19[53],x_20[53],x_21[53],x_22[53],x_23[53],x_24[53],x_25[53],x_26[53],x_27[53],x_28[53],x_29[53],x_30[53],x_31[53],x_32[53]}),.c_in(c_in_53),.c_out(c_in_54),.s(s_53),.c(c_53));
wire  c_54;
wire  s_54;
wallace_tree_ w54(.clk(clk),.rst_n(rst_n),.a({x_0[54],x_1[54],x_2[54],x_3[54],x_4[54],x_5[54],x_6[54],x_7[54],x_8[54],x_9[54],x_10[54],x_11[54],x_12[54],x_13[54],x_14[54],x_15[54],x_16[54],x_17[54],x_18[54],x_19[54],x_20[54],x_21[54],x_22[54],x_23[54],x_24[54],x_25[54],x_26[54],x_27[54],x_28[54],x_29[54],x_30[54],x_31[54],x_32[54]}),.c_in(c_in_54),.c_out(c_in_55),.s(s_54),.c(c_54));
wire  c_55;
wire  s_55;
wallace_tree_ w55(.clk(clk),.rst_n(rst_n),.a({x_0[55],x_1[55],x_2[55],x_3[55],x_4[55],x_5[55],x_6[55],x_7[55],x_8[55],x_9[55],x_10[55],x_11[55],x_12[55],x_13[55],x_14[55],x_15[55],x_16[55],x_17[55],x_18[55],x_19[55],x_20[55],x_21[55],x_22[55],x_23[55],x_24[55],x_25[55],x_26[55],x_27[55],x_28[55],x_29[55],x_30[55],x_31[55],x_32[55]}),.c_in(c_in_55),.c_out(c_in_56),.s(s_55),.c(c_55));
wire  c_56;
wire  s_56;
wallace_tree_ w56(.clk(clk),.rst_n(rst_n),.a({x_0[56],x_1[56],x_2[56],x_3[56],x_4[56],x_5[56],x_6[56],x_7[56],x_8[56],x_9[56],x_10[56],x_11[56],x_12[56],x_13[56],x_14[56],x_15[56],x_16[56],x_17[56],x_18[56],x_19[56],x_20[56],x_21[56],x_22[56],x_23[56],x_24[56],x_25[56],x_26[56],x_27[56],x_28[56],x_29[56],x_30[56],x_31[56],x_32[56]}),.c_in(c_in_56),.c_out(c_in_57),.s(s_56),.c(c_56));
wire  c_57;
wire  s_57;
wallace_tree_ w57(.clk(clk),.rst_n(rst_n),.a({x_0[57],x_1[57],x_2[57],x_3[57],x_4[57],x_5[57],x_6[57],x_7[57],x_8[57],x_9[57],x_10[57],x_11[57],x_12[57],x_13[57],x_14[57],x_15[57],x_16[57],x_17[57],x_18[57],x_19[57],x_20[57],x_21[57],x_22[57],x_23[57],x_24[57],x_25[57],x_26[57],x_27[57],x_28[57],x_29[57],x_30[57],x_31[57],x_32[57]}),.c_in(c_in_57),.c_out(c_in_58),.s(s_57),.c(c_57));
wire  c_58;
wire  s_58;
wallace_tree_ w58(.clk(clk),.rst_n(rst_n),.a({x_0[58],x_1[58],x_2[58],x_3[58],x_4[58],x_5[58],x_6[58],x_7[58],x_8[58],x_9[58],x_10[58],x_11[58],x_12[58],x_13[58],x_14[58],x_15[58],x_16[58],x_17[58],x_18[58],x_19[58],x_20[58],x_21[58],x_22[58],x_23[58],x_24[58],x_25[58],x_26[58],x_27[58],x_28[58],x_29[58],x_30[58],x_31[58],x_32[58]}),.c_in(c_in_58),.c_out(c_in_59),.s(s_58),.c(c_58));
wire  c_59;
wire  s_59;
wallace_tree_ w59(.clk(clk),.rst_n(rst_n),.a({x_0[59],x_1[59],x_2[59],x_3[59],x_4[59],x_5[59],x_6[59],x_7[59],x_8[59],x_9[59],x_10[59],x_11[59],x_12[59],x_13[59],x_14[59],x_15[59],x_16[59],x_17[59],x_18[59],x_19[59],x_20[59],x_21[59],x_22[59],x_23[59],x_24[59],x_25[59],x_26[59],x_27[59],x_28[59],x_29[59],x_30[59],x_31[59],x_32[59]}),.c_in(c_in_59),.c_out(c_in_60),.s(s_59),.c(c_59));
wire  c_60;
wire  s_60;
wallace_tree_ w60(.clk(clk),.rst_n(rst_n),.a({x_0[60],x_1[60],x_2[60],x_3[60],x_4[60],x_5[60],x_6[60],x_7[60],x_8[60],x_9[60],x_10[60],x_11[60],x_12[60],x_13[60],x_14[60],x_15[60],x_16[60],x_17[60],x_18[60],x_19[60],x_20[60],x_21[60],x_22[60],x_23[60],x_24[60],x_25[60],x_26[60],x_27[60],x_28[60],x_29[60],x_30[60],x_31[60],x_32[60]}),.c_in(c_in_60),.c_out(c_in_61),.s(s_60),.c(c_60));
wire  c_61;
wire  s_61;
wallace_tree_ w61(.clk(clk),.rst_n(rst_n),.a({x_0[61],x_1[61],x_2[61],x_3[61],x_4[61],x_5[61],x_6[61],x_7[61],x_8[61],x_9[61],x_10[61],x_11[61],x_12[61],x_13[61],x_14[61],x_15[61],x_16[61],x_17[61],x_18[61],x_19[61],x_20[61],x_21[61],x_22[61],x_23[61],x_24[61],x_25[61],x_26[61],x_27[61],x_28[61],x_29[61],x_30[61],x_31[61],x_32[61]}),.c_in(c_in_61),.c_out(c_in_62),.s(s_61),.c(c_61));
wire  c_62;
wire  s_62;
wallace_tree_ w62(.clk(clk),.rst_n(rst_n),.a({x_0[62],x_1[62],x_2[62],x_3[62],x_4[62],x_5[62],x_6[62],x_7[62],x_8[62],x_9[62],x_10[62],x_11[62],x_12[62],x_13[62],x_14[62],x_15[62],x_16[62],x_17[62],x_18[62],x_19[62],x_20[62],x_21[62],x_22[62],x_23[62],x_24[62],x_25[62],x_26[62],x_27[62],x_28[62],x_29[62],x_30[62],x_31[62],x_32[62]}),.c_in(c_in_62),.c_out(c_in_63),.s(s_62),.c(c_62));
wire  c_63;
wire  s_63;
wallace_tree_ w63(.clk(clk),.rst_n(rst_n),.a({x_0[63],x_1[63],x_2[63],x_3[63],x_4[63],x_5[63],x_6[63],x_7[63],x_8[63],x_9[63],x_10[63],x_11[63],x_12[63],x_13[63],x_14[63],x_15[63],x_16[63],x_17[63],x_18[63],x_19[63],x_20[63],x_21[63],x_22[63],x_23[63],x_24[63],x_25[63],x_26[63],x_27[63],x_28[63],x_29[63],x_30[63],x_31[63],x_32[63]}),.c_in(c_in_63),.c_out(c_in_64),.s(s_63),.c(c_63));
wire  c_64;
wire  s_64;
wallace_tree_ w64(.clk(clk),.rst_n(rst_n),.a({x_0[64],x_1[64],x_2[64],x_3[64],x_4[64],x_5[64],x_6[64],x_7[64],x_8[64],x_9[64],x_10[64],x_11[64],x_12[64],x_13[64],x_14[64],x_15[64],x_16[64],x_17[64],x_18[64],x_19[64],x_20[64],x_21[64],x_22[64],x_23[64],x_24[64],x_25[64],x_26[64],x_27[64],x_28[64],x_29[64],x_30[64],x_31[64],x_32[64]}),.c_in(c_in_64),.c_out(c_in_65),.s(s_64),.c(c_64));
wire  c_65;
wire  s_65;
wallace_tree_ w65(.clk(clk),.rst_n(rst_n),.a({x_0[65],x_1[65],x_2[65],x_3[65],x_4[65],x_5[65],x_6[65],x_7[65],x_8[65],x_9[65],x_10[65],x_11[65],x_12[65],x_13[65],x_14[65],x_15[65],x_16[65],x_17[65],x_18[65],x_19[65],x_20[65],x_21[65],x_22[65],x_23[65],x_24[65],x_25[65],x_26[65],x_27[65],x_28[65],x_29[65],x_30[65],x_31[65],x_32[65]}),.c_in(c_in_65),.c_out(c_in_66),.s(s_65),.c(c_65));
wire  c_66;
wire  s_66;
wallace_tree_ w66(.clk(clk),.rst_n(rst_n),.a({x_0[66],x_1[66],x_2[66],x_3[66],x_4[66],x_5[66],x_6[66],x_7[66],x_8[66],x_9[66],x_10[66],x_11[66],x_12[66],x_13[66],x_14[66],x_15[66],x_16[66],x_17[66],x_18[66],x_19[66],x_20[66],x_21[66],x_22[66],x_23[66],x_24[66],x_25[66],x_26[66],x_27[66],x_28[66],x_29[66],x_30[66],x_31[66],x_32[66]}),.c_in(c_in_66),.c_out(c_in_67),.s(s_66),.c(c_66));
wire  c_67;
wire  s_67;
wallace_tree_ w67(.clk(clk),.rst_n(rst_n),.a({x_0[67],x_1[67],x_2[67],x_3[67],x_4[67],x_5[67],x_6[67],x_7[67],x_8[67],x_9[67],x_10[67],x_11[67],x_12[67],x_13[67],x_14[67],x_15[67],x_16[67],x_17[67],x_18[67],x_19[67],x_20[67],x_21[67],x_22[67],x_23[67],x_24[67],x_25[67],x_26[67],x_27[67],x_28[67],x_29[67],x_30[67],x_31[67],x_32[67]}),.c_in(c_in_67),.c_out(c_in_68),.s(s_67),.c(c_67));
wire  c_68;
wire  s_68;
wallace_tree_ w68(.clk(clk),.rst_n(rst_n),.a({x_0[68],x_1[68],x_2[68],x_3[68],x_4[68],x_5[68],x_6[68],x_7[68],x_8[68],x_9[68],x_10[68],x_11[68],x_12[68],x_13[68],x_14[68],x_15[68],x_16[68],x_17[68],x_18[68],x_19[68],x_20[68],x_21[68],x_22[68],x_23[68],x_24[68],x_25[68],x_26[68],x_27[68],x_28[68],x_29[68],x_30[68],x_31[68],x_32[68]}),.c_in(c_in_68),.c_out(c_in_69),.s(s_68),.c(c_68));
wire  c_69;
wire  s_69;
wallace_tree_ w69(.clk(clk),.rst_n(rst_n),.a({x_0[69],x_1[69],x_2[69],x_3[69],x_4[69],x_5[69],x_6[69],x_7[69],x_8[69],x_9[69],x_10[69],x_11[69],x_12[69],x_13[69],x_14[69],x_15[69],x_16[69],x_17[69],x_18[69],x_19[69],x_20[69],x_21[69],x_22[69],x_23[69],x_24[69],x_25[69],x_26[69],x_27[69],x_28[69],x_29[69],x_30[69],x_31[69],x_32[69]}),.c_in(c_in_69),.c_out(c_in_70),.s(s_69),.c(c_69));
wire  c_70;
wire  s_70;
wallace_tree_ w70(.clk(clk),.rst_n(rst_n),.a({x_0[70],x_1[70],x_2[70],x_3[70],x_4[70],x_5[70],x_6[70],x_7[70],x_8[70],x_9[70],x_10[70],x_11[70],x_12[70],x_13[70],x_14[70],x_15[70],x_16[70],x_17[70],x_18[70],x_19[70],x_20[70],x_21[70],x_22[70],x_23[70],x_24[70],x_25[70],x_26[70],x_27[70],x_28[70],x_29[70],x_30[70],x_31[70],x_32[70]}),.c_in(c_in_70),.c_out(c_in_71),.s(s_70),.c(c_70));
wire  c_71;
wire  s_71;
wallace_tree_ w71(.clk(clk),.rst_n(rst_n),.a({x_0[71],x_1[71],x_2[71],x_3[71],x_4[71],x_5[71],x_6[71],x_7[71],x_8[71],x_9[71],x_10[71],x_11[71],x_12[71],x_13[71],x_14[71],x_15[71],x_16[71],x_17[71],x_18[71],x_19[71],x_20[71],x_21[71],x_22[71],x_23[71],x_24[71],x_25[71],x_26[71],x_27[71],x_28[71],x_29[71],x_30[71],x_31[71],x_32[71]}),.c_in(c_in_71),.c_out(c_in_72),.s(s_71),.c(c_71));
wire  c_72;
wire  s_72;
wallace_tree_ w72(.clk(clk),.rst_n(rst_n),.a({x_0[72],x_1[72],x_2[72],x_3[72],x_4[72],x_5[72],x_6[72],x_7[72],x_8[72],x_9[72],x_10[72],x_11[72],x_12[72],x_13[72],x_14[72],x_15[72],x_16[72],x_17[72],x_18[72],x_19[72],x_20[72],x_21[72],x_22[72],x_23[72],x_24[72],x_25[72],x_26[72],x_27[72],x_28[72],x_29[72],x_30[72],x_31[72],x_32[72]}),.c_in(c_in_72),.c_out(c_in_73),.s(s_72),.c(c_72));
wire  c_73;
wire  s_73;
wallace_tree_ w73(.clk(clk),.rst_n(rst_n),.a({x_0[73],x_1[73],x_2[73],x_3[73],x_4[73],x_5[73],x_6[73],x_7[73],x_8[73],x_9[73],x_10[73],x_11[73],x_12[73],x_13[73],x_14[73],x_15[73],x_16[73],x_17[73],x_18[73],x_19[73],x_20[73],x_21[73],x_22[73],x_23[73],x_24[73],x_25[73],x_26[73],x_27[73],x_28[73],x_29[73],x_30[73],x_31[73],x_32[73]}),.c_in(c_in_73),.c_out(c_in_74),.s(s_73),.c(c_73));
wire  c_74;
wire  s_74;
wallace_tree_ w74(.clk(clk),.rst_n(rst_n),.a({x_0[74],x_1[74],x_2[74],x_3[74],x_4[74],x_5[74],x_6[74],x_7[74],x_8[74],x_9[74],x_10[74],x_11[74],x_12[74],x_13[74],x_14[74],x_15[74],x_16[74],x_17[74],x_18[74],x_19[74],x_20[74],x_21[74],x_22[74],x_23[74],x_24[74],x_25[74],x_26[74],x_27[74],x_28[74],x_29[74],x_30[74],x_31[74],x_32[74]}),.c_in(c_in_74),.c_out(c_in_75),.s(s_74),.c(c_74));
wire  c_75;
wire  s_75;
wallace_tree_ w75(.clk(clk),.rst_n(rst_n),.a({x_0[75],x_1[75],x_2[75],x_3[75],x_4[75],x_5[75],x_6[75],x_7[75],x_8[75],x_9[75],x_10[75],x_11[75],x_12[75],x_13[75],x_14[75],x_15[75],x_16[75],x_17[75],x_18[75],x_19[75],x_20[75],x_21[75],x_22[75],x_23[75],x_24[75],x_25[75],x_26[75],x_27[75],x_28[75],x_29[75],x_30[75],x_31[75],x_32[75]}),.c_in(c_in_75),.c_out(c_in_76),.s(s_75),.c(c_75));
wire  c_76;
wire  s_76;
wallace_tree_ w76(.clk(clk),.rst_n(rst_n),.a({x_0[76],x_1[76],x_2[76],x_3[76],x_4[76],x_5[76],x_6[76],x_7[76],x_8[76],x_9[76],x_10[76],x_11[76],x_12[76],x_13[76],x_14[76],x_15[76],x_16[76],x_17[76],x_18[76],x_19[76],x_20[76],x_21[76],x_22[76],x_23[76],x_24[76],x_25[76],x_26[76],x_27[76],x_28[76],x_29[76],x_30[76],x_31[76],x_32[76]}),.c_in(c_in_76),.c_out(c_in_77),.s(s_76),.c(c_76));
wire  c_77;
wire  s_77;
wallace_tree_ w77(.clk(clk),.rst_n(rst_n),.a({x_0[77],x_1[77],x_2[77],x_3[77],x_4[77],x_5[77],x_6[77],x_7[77],x_8[77],x_9[77],x_10[77],x_11[77],x_12[77],x_13[77],x_14[77],x_15[77],x_16[77],x_17[77],x_18[77],x_19[77],x_20[77],x_21[77],x_22[77],x_23[77],x_24[77],x_25[77],x_26[77],x_27[77],x_28[77],x_29[77],x_30[77],x_31[77],x_32[77]}),.c_in(c_in_77),.c_out(c_in_78),.s(s_77),.c(c_77));
wire  c_78;
wire  s_78;
wallace_tree_ w78(.clk(clk),.rst_n(rst_n),.a({x_0[78],x_1[78],x_2[78],x_3[78],x_4[78],x_5[78],x_6[78],x_7[78],x_8[78],x_9[78],x_10[78],x_11[78],x_12[78],x_13[78],x_14[78],x_15[78],x_16[78],x_17[78],x_18[78],x_19[78],x_20[78],x_21[78],x_22[78],x_23[78],x_24[78],x_25[78],x_26[78],x_27[78],x_28[78],x_29[78],x_30[78],x_31[78],x_32[78]}),.c_in(c_in_78),.c_out(c_in_79),.s(s_78),.c(c_78));
wire  c_79;
wire  s_79;
wallace_tree_ w79(.clk(clk),.rst_n(rst_n),.a({x_0[79],x_1[79],x_2[79],x_3[79],x_4[79],x_5[79],x_6[79],x_7[79],x_8[79],x_9[79],x_10[79],x_11[79],x_12[79],x_13[79],x_14[79],x_15[79],x_16[79],x_17[79],x_18[79],x_19[79],x_20[79],x_21[79],x_22[79],x_23[79],x_24[79],x_25[79],x_26[79],x_27[79],x_28[79],x_29[79],x_30[79],x_31[79],x_32[79]}),.c_in(c_in_79),.c_out(c_in_80),.s(s_79),.c(c_79));
wire  c_80;
wire  s_80;
wallace_tree_ w80(.clk(clk),.rst_n(rst_n),.a({x_0[80],x_1[80],x_2[80],x_3[80],x_4[80],x_5[80],x_6[80],x_7[80],x_8[80],x_9[80],x_10[80],x_11[80],x_12[80],x_13[80],x_14[80],x_15[80],x_16[80],x_17[80],x_18[80],x_19[80],x_20[80],x_21[80],x_22[80],x_23[80],x_24[80],x_25[80],x_26[80],x_27[80],x_28[80],x_29[80],x_30[80],x_31[80],x_32[80]}),.c_in(c_in_80),.c_out(c_in_81),.s(s_80),.c(c_80));
wire  c_81;
wire  s_81;
wallace_tree_ w81(.clk(clk),.rst_n(rst_n),.a({x_0[81],x_1[81],x_2[81],x_3[81],x_4[81],x_5[81],x_6[81],x_7[81],x_8[81],x_9[81],x_10[81],x_11[81],x_12[81],x_13[81],x_14[81],x_15[81],x_16[81],x_17[81],x_18[81],x_19[81],x_20[81],x_21[81],x_22[81],x_23[81],x_24[81],x_25[81],x_26[81],x_27[81],x_28[81],x_29[81],x_30[81],x_31[81],x_32[81]}),.c_in(c_in_81),.c_out(c_in_82),.s(s_81),.c(c_81));
wire  c_82;
wire  s_82;
wallace_tree_ w82(.clk(clk),.rst_n(rst_n),.a({x_0[82],x_1[82],x_2[82],x_3[82],x_4[82],x_5[82],x_6[82],x_7[82],x_8[82],x_9[82],x_10[82],x_11[82],x_12[82],x_13[82],x_14[82],x_15[82],x_16[82],x_17[82],x_18[82],x_19[82],x_20[82],x_21[82],x_22[82],x_23[82],x_24[82],x_25[82],x_26[82],x_27[82],x_28[82],x_29[82],x_30[82],x_31[82],x_32[82]}),.c_in(c_in_82),.c_out(c_in_83),.s(s_82),.c(c_82));
wire  c_83;
wire  s_83;
wallace_tree_ w83(.clk(clk),.rst_n(rst_n),.a({x_0[83],x_1[83],x_2[83],x_3[83],x_4[83],x_5[83],x_6[83],x_7[83],x_8[83],x_9[83],x_10[83],x_11[83],x_12[83],x_13[83],x_14[83],x_15[83],x_16[83],x_17[83],x_18[83],x_19[83],x_20[83],x_21[83],x_22[83],x_23[83],x_24[83],x_25[83],x_26[83],x_27[83],x_28[83],x_29[83],x_30[83],x_31[83],x_32[83]}),.c_in(c_in_83),.c_out(c_in_84),.s(s_83),.c(c_83));
wire  c_84;
wire  s_84;
wallace_tree_ w84(.clk(clk),.rst_n(rst_n),.a({x_0[84],x_1[84],x_2[84],x_3[84],x_4[84],x_5[84],x_6[84],x_7[84],x_8[84],x_9[84],x_10[84],x_11[84],x_12[84],x_13[84],x_14[84],x_15[84],x_16[84],x_17[84],x_18[84],x_19[84],x_20[84],x_21[84],x_22[84],x_23[84],x_24[84],x_25[84],x_26[84],x_27[84],x_28[84],x_29[84],x_30[84],x_31[84],x_32[84]}),.c_in(c_in_84),.c_out(c_in_85),.s(s_84),.c(c_84));
wire  c_85;
wire  s_85;
wallace_tree_ w85(.clk(clk),.rst_n(rst_n),.a({x_0[85],x_1[85],x_2[85],x_3[85],x_4[85],x_5[85],x_6[85],x_7[85],x_8[85],x_9[85],x_10[85],x_11[85],x_12[85],x_13[85],x_14[85],x_15[85],x_16[85],x_17[85],x_18[85],x_19[85],x_20[85],x_21[85],x_22[85],x_23[85],x_24[85],x_25[85],x_26[85],x_27[85],x_28[85],x_29[85],x_30[85],x_31[85],x_32[85]}),.c_in(c_in_85),.c_out(c_in_86),.s(s_85),.c(c_85));
wire  c_86;
wire  s_86;
wallace_tree_ w86(.clk(clk),.rst_n(rst_n),.a({x_0[86],x_1[86],x_2[86],x_3[86],x_4[86],x_5[86],x_6[86],x_7[86],x_8[86],x_9[86],x_10[86],x_11[86],x_12[86],x_13[86],x_14[86],x_15[86],x_16[86],x_17[86],x_18[86],x_19[86],x_20[86],x_21[86],x_22[86],x_23[86],x_24[86],x_25[86],x_26[86],x_27[86],x_28[86],x_29[86],x_30[86],x_31[86],x_32[86]}),.c_in(c_in_86),.c_out(c_in_87),.s(s_86),.c(c_86));
wire  c_87;
wire  s_87;
wallace_tree_ w87(.clk(clk),.rst_n(rst_n),.a({x_0[87],x_1[87],x_2[87],x_3[87],x_4[87],x_5[87],x_6[87],x_7[87],x_8[87],x_9[87],x_10[87],x_11[87],x_12[87],x_13[87],x_14[87],x_15[87],x_16[87],x_17[87],x_18[87],x_19[87],x_20[87],x_21[87],x_22[87],x_23[87],x_24[87],x_25[87],x_26[87],x_27[87],x_28[87],x_29[87],x_30[87],x_31[87],x_32[87]}),.c_in(c_in_87),.c_out(c_in_88),.s(s_87),.c(c_87));
wire  c_88;
wire  s_88;
wallace_tree_ w88(.clk(clk),.rst_n(rst_n),.a({x_0[88],x_1[88],x_2[88],x_3[88],x_4[88],x_5[88],x_6[88],x_7[88],x_8[88],x_9[88],x_10[88],x_11[88],x_12[88],x_13[88],x_14[88],x_15[88],x_16[88],x_17[88],x_18[88],x_19[88],x_20[88],x_21[88],x_22[88],x_23[88],x_24[88],x_25[88],x_26[88],x_27[88],x_28[88],x_29[88],x_30[88],x_31[88],x_32[88]}),.c_in(c_in_88),.c_out(c_in_89),.s(s_88),.c(c_88));
wire  c_89;
wire  s_89;
wallace_tree_ w89(.clk(clk),.rst_n(rst_n),.a({x_0[89],x_1[89],x_2[89],x_3[89],x_4[89],x_5[89],x_6[89],x_7[89],x_8[89],x_9[89],x_10[89],x_11[89],x_12[89],x_13[89],x_14[89],x_15[89],x_16[89],x_17[89],x_18[89],x_19[89],x_20[89],x_21[89],x_22[89],x_23[89],x_24[89],x_25[89],x_26[89],x_27[89],x_28[89],x_29[89],x_30[89],x_31[89],x_32[89]}),.c_in(c_in_89),.c_out(c_in_90),.s(s_89),.c(c_89));
wire  c_90;
wire  s_90;
wallace_tree_ w90(.clk(clk),.rst_n(rst_n),.a({x_0[90],x_1[90],x_2[90],x_3[90],x_4[90],x_5[90],x_6[90],x_7[90],x_8[90],x_9[90],x_10[90],x_11[90],x_12[90],x_13[90],x_14[90],x_15[90],x_16[90],x_17[90],x_18[90],x_19[90],x_20[90],x_21[90],x_22[90],x_23[90],x_24[90],x_25[90],x_26[90],x_27[90],x_28[90],x_29[90],x_30[90],x_31[90],x_32[90]}),.c_in(c_in_90),.c_out(c_in_91),.s(s_90),.c(c_90));
wire  c_91;
wire  s_91;
wallace_tree_ w91(.clk(clk),.rst_n(rst_n),.a({x_0[91],x_1[91],x_2[91],x_3[91],x_4[91],x_5[91],x_6[91],x_7[91],x_8[91],x_9[91],x_10[91],x_11[91],x_12[91],x_13[91],x_14[91],x_15[91],x_16[91],x_17[91],x_18[91],x_19[91],x_20[91],x_21[91],x_22[91],x_23[91],x_24[91],x_25[91],x_26[91],x_27[91],x_28[91],x_29[91],x_30[91],x_31[91],x_32[91]}),.c_in(c_in_91),.c_out(c_in_92),.s(s_91),.c(c_91));
wire  c_92;
wire  s_92;
wallace_tree_ w92(.clk(clk),.rst_n(rst_n),.a({x_0[92],x_1[92],x_2[92],x_3[92],x_4[92],x_5[92],x_6[92],x_7[92],x_8[92],x_9[92],x_10[92],x_11[92],x_12[92],x_13[92],x_14[92],x_15[92],x_16[92],x_17[92],x_18[92],x_19[92],x_20[92],x_21[92],x_22[92],x_23[92],x_24[92],x_25[92],x_26[92],x_27[92],x_28[92],x_29[92],x_30[92],x_31[92],x_32[92]}),.c_in(c_in_92),.c_out(c_in_93),.s(s_92),.c(c_92));
wire  c_93;
wire  s_93;
wallace_tree_ w93(.clk(clk),.rst_n(rst_n),.a({x_0[93],x_1[93],x_2[93],x_3[93],x_4[93],x_5[93],x_6[93],x_7[93],x_8[93],x_9[93],x_10[93],x_11[93],x_12[93],x_13[93],x_14[93],x_15[93],x_16[93],x_17[93],x_18[93],x_19[93],x_20[93],x_21[93],x_22[93],x_23[93],x_24[93],x_25[93],x_26[93],x_27[93],x_28[93],x_29[93],x_30[93],x_31[93],x_32[93]}),.c_in(c_in_93),.c_out(c_in_94),.s(s_93),.c(c_93));
wire  c_94;
wire  s_94;
wallace_tree_ w94(.clk(clk),.rst_n(rst_n),.a({x_0[94],x_1[94],x_2[94],x_3[94],x_4[94],x_5[94],x_6[94],x_7[94],x_8[94],x_9[94],x_10[94],x_11[94],x_12[94],x_13[94],x_14[94],x_15[94],x_16[94],x_17[94],x_18[94],x_19[94],x_20[94],x_21[94],x_22[94],x_23[94],x_24[94],x_25[94],x_26[94],x_27[94],x_28[94],x_29[94],x_30[94],x_31[94],x_32[94]}),.c_in(c_in_94),.c_out(c_in_95),.s(s_94),.c(c_94));
wire  c_95;
wire  s_95;
wallace_tree_ w95(.clk(clk),.rst_n(rst_n),.a({x_0[95],x_1[95],x_2[95],x_3[95],x_4[95],x_5[95],x_6[95],x_7[95],x_8[95],x_9[95],x_10[95],x_11[95],x_12[95],x_13[95],x_14[95],x_15[95],x_16[95],x_17[95],x_18[95],x_19[95],x_20[95],x_21[95],x_22[95],x_23[95],x_24[95],x_25[95],x_26[95],x_27[95],x_28[95],x_29[95],x_30[95],x_31[95],x_32[95]}),.c_in(c_in_95),.c_out(c_in_96),.s(s_95),.c(c_95));
wire  c_96;
wire  s_96;
wallace_tree_ w96(.clk(clk),.rst_n(rst_n),.a({x_0[96],x_1[96],x_2[96],x_3[96],x_4[96],x_5[96],x_6[96],x_7[96],x_8[96],x_9[96],x_10[96],x_11[96],x_12[96],x_13[96],x_14[96],x_15[96],x_16[96],x_17[96],x_18[96],x_19[96],x_20[96],x_21[96],x_22[96],x_23[96],x_24[96],x_25[96],x_26[96],x_27[96],x_28[96],x_29[96],x_30[96],x_31[96],x_32[96]}),.c_in(c_in_96),.c_out(c_in_97),.s(s_96),.c(c_96));
wire  c_97;
wire  s_97;
wallace_tree_ w97(.clk(clk),.rst_n(rst_n),.a({x_0[97],x_1[97],x_2[97],x_3[97],x_4[97],x_5[97],x_6[97],x_7[97],x_8[97],x_9[97],x_10[97],x_11[97],x_12[97],x_13[97],x_14[97],x_15[97],x_16[97],x_17[97],x_18[97],x_19[97],x_20[97],x_21[97],x_22[97],x_23[97],x_24[97],x_25[97],x_26[97],x_27[97],x_28[97],x_29[97],x_30[97],x_31[97],x_32[97]}),.c_in(c_in_97),.c_out(c_in_98),.s(s_97),.c(c_97));
wire  c_98;
wire  s_98;
wallace_tree_ w98(.clk(clk),.rst_n(rst_n),.a({x_0[98],x_1[98],x_2[98],x_3[98],x_4[98],x_5[98],x_6[98],x_7[98],x_8[98],x_9[98],x_10[98],x_11[98],x_12[98],x_13[98],x_14[98],x_15[98],x_16[98],x_17[98],x_18[98],x_19[98],x_20[98],x_21[98],x_22[98],x_23[98],x_24[98],x_25[98],x_26[98],x_27[98],x_28[98],x_29[98],x_30[98],x_31[98],x_32[98]}),.c_in(c_in_98),.c_out(c_in_99),.s(s_98),.c(c_98));
wire  c_99;
wire  s_99;
wallace_tree_ w99(.clk(clk),.rst_n(rst_n),.a({x_0[99],x_1[99],x_2[99],x_3[99],x_4[99],x_5[99],x_6[99],x_7[99],x_8[99],x_9[99],x_10[99],x_11[99],x_12[99],x_13[99],x_14[99],x_15[99],x_16[99],x_17[99],x_18[99],x_19[99],x_20[99],x_21[99],x_22[99],x_23[99],x_24[99],x_25[99],x_26[99],x_27[99],x_28[99],x_29[99],x_30[99],x_31[99],x_32[99]}),.c_in(c_in_99),.c_out(c_in_100),.s(s_99),.c(c_99));
wire  c_100;
wire  s_100;
wallace_tree_ w100(.clk(clk),.rst_n(rst_n),.a({x_0[100],x_1[100],x_2[100],x_3[100],x_4[100],x_5[100],x_6[100],x_7[100],x_8[100],x_9[100],x_10[100],x_11[100],x_12[100],x_13[100],x_14[100],x_15[100],x_16[100],x_17[100],x_18[100],x_19[100],x_20[100],x_21[100],x_22[100],x_23[100],x_24[100],x_25[100],x_26[100],x_27[100],x_28[100],x_29[100],x_30[100],x_31[100],x_32[100]}),.c_in(c_in_100),.c_out(c_in_101),.s(s_100),.c(c_100));
wire  c_101;
wire  s_101;
wallace_tree_ w101(.clk(clk),.rst_n(rst_n),.a({x_0[101],x_1[101],x_2[101],x_3[101],x_4[101],x_5[101],x_6[101],x_7[101],x_8[101],x_9[101],x_10[101],x_11[101],x_12[101],x_13[101],x_14[101],x_15[101],x_16[101],x_17[101],x_18[101],x_19[101],x_20[101],x_21[101],x_22[101],x_23[101],x_24[101],x_25[101],x_26[101],x_27[101],x_28[101],x_29[101],x_30[101],x_31[101],x_32[101]}),.c_in(c_in_101),.c_out(c_in_102),.s(s_101),.c(c_101));
wire  c_102;
wire  s_102;
wallace_tree_ w102(.clk(clk),.rst_n(rst_n),.a({x_0[102],x_1[102],x_2[102],x_3[102],x_4[102],x_5[102],x_6[102],x_7[102],x_8[102],x_9[102],x_10[102],x_11[102],x_12[102],x_13[102],x_14[102],x_15[102],x_16[102],x_17[102],x_18[102],x_19[102],x_20[102],x_21[102],x_22[102],x_23[102],x_24[102],x_25[102],x_26[102],x_27[102],x_28[102],x_29[102],x_30[102],x_31[102],x_32[102]}),.c_in(c_in_102),.c_out(c_in_103),.s(s_102),.c(c_102));
wire  c_103;
wire  s_103;
wallace_tree_ w103(.clk(clk),.rst_n(rst_n),.a({x_0[103],x_1[103],x_2[103],x_3[103],x_4[103],x_5[103],x_6[103],x_7[103],x_8[103],x_9[103],x_10[103],x_11[103],x_12[103],x_13[103],x_14[103],x_15[103],x_16[103],x_17[103],x_18[103],x_19[103],x_20[103],x_21[103],x_22[103],x_23[103],x_24[103],x_25[103],x_26[103],x_27[103],x_28[103],x_29[103],x_30[103],x_31[103],x_32[103]}),.c_in(c_in_103),.c_out(c_in_104),.s(s_103),.c(c_103));
wire  c_104;
wire  s_104;
wallace_tree_ w104(.clk(clk),.rst_n(rst_n),.a({x_0[104],x_1[104],x_2[104],x_3[104],x_4[104],x_5[104],x_6[104],x_7[104],x_8[104],x_9[104],x_10[104],x_11[104],x_12[104],x_13[104],x_14[104],x_15[104],x_16[104],x_17[104],x_18[104],x_19[104],x_20[104],x_21[104],x_22[104],x_23[104],x_24[104],x_25[104],x_26[104],x_27[104],x_28[104],x_29[104],x_30[104],x_31[104],x_32[104]}),.c_in(c_in_104),.c_out(c_in_105),.s(s_104),.c(c_104));
wire  c_105;
wire  s_105;
wallace_tree_ w105(.clk(clk),.rst_n(rst_n),.a({x_0[105],x_1[105],x_2[105],x_3[105],x_4[105],x_5[105],x_6[105],x_7[105],x_8[105],x_9[105],x_10[105],x_11[105],x_12[105],x_13[105],x_14[105],x_15[105],x_16[105],x_17[105],x_18[105],x_19[105],x_20[105],x_21[105],x_22[105],x_23[105],x_24[105],x_25[105],x_26[105],x_27[105],x_28[105],x_29[105],x_30[105],x_31[105],x_32[105]}),.c_in(c_in_105),.c_out(c_in_106),.s(s_105),.c(c_105));
wire  c_106;
wire  s_106;
wallace_tree_ w106(.clk(clk),.rst_n(rst_n),.a({x_0[106],x_1[106],x_2[106],x_3[106],x_4[106],x_5[106],x_6[106],x_7[106],x_8[106],x_9[106],x_10[106],x_11[106],x_12[106],x_13[106],x_14[106],x_15[106],x_16[106],x_17[106],x_18[106],x_19[106],x_20[106],x_21[106],x_22[106],x_23[106],x_24[106],x_25[106],x_26[106],x_27[106],x_28[106],x_29[106],x_30[106],x_31[106],x_32[106]}),.c_in(c_in_106),.c_out(c_in_107),.s(s_106),.c(c_106));
wire  c_107;
wire  s_107;
wallace_tree_ w107(.clk(clk),.rst_n(rst_n),.a({x_0[107],x_1[107],x_2[107],x_3[107],x_4[107],x_5[107],x_6[107],x_7[107],x_8[107],x_9[107],x_10[107],x_11[107],x_12[107],x_13[107],x_14[107],x_15[107],x_16[107],x_17[107],x_18[107],x_19[107],x_20[107],x_21[107],x_22[107],x_23[107],x_24[107],x_25[107],x_26[107],x_27[107],x_28[107],x_29[107],x_30[107],x_31[107],x_32[107]}),.c_in(c_in_107),.c_out(c_in_108),.s(s_107),.c(c_107));
wire  c_108;
wire  s_108;
wallace_tree_ w108(.clk(clk),.rst_n(rst_n),.a({x_0[108],x_1[108],x_2[108],x_3[108],x_4[108],x_5[108],x_6[108],x_7[108],x_8[108],x_9[108],x_10[108],x_11[108],x_12[108],x_13[108],x_14[108],x_15[108],x_16[108],x_17[108],x_18[108],x_19[108],x_20[108],x_21[108],x_22[108],x_23[108],x_24[108],x_25[108],x_26[108],x_27[108],x_28[108],x_29[108],x_30[108],x_31[108],x_32[108]}),.c_in(c_in_108),.c_out(c_in_109),.s(s_108),.c(c_108));
wire  c_109;
wire  s_109;
wallace_tree_ w109(.clk(clk),.rst_n(rst_n),.a({x_0[109],x_1[109],x_2[109],x_3[109],x_4[109],x_5[109],x_6[109],x_7[109],x_8[109],x_9[109],x_10[109],x_11[109],x_12[109],x_13[109],x_14[109],x_15[109],x_16[109],x_17[109],x_18[109],x_19[109],x_20[109],x_21[109],x_22[109],x_23[109],x_24[109],x_25[109],x_26[109],x_27[109],x_28[109],x_29[109],x_30[109],x_31[109],x_32[109]}),.c_in(c_in_109),.c_out(c_in_110),.s(s_109),.c(c_109));
wire  c_110;
wire  s_110;
wallace_tree_ w110(.clk(clk),.rst_n(rst_n),.a({x_0[110],x_1[110],x_2[110],x_3[110],x_4[110],x_5[110],x_6[110],x_7[110],x_8[110],x_9[110],x_10[110],x_11[110],x_12[110],x_13[110],x_14[110],x_15[110],x_16[110],x_17[110],x_18[110],x_19[110],x_20[110],x_21[110],x_22[110],x_23[110],x_24[110],x_25[110],x_26[110],x_27[110],x_28[110],x_29[110],x_30[110],x_31[110],x_32[110]}),.c_in(c_in_110),.c_out(c_in_111),.s(s_110),.c(c_110));
wire  c_111;
wire  s_111;
wallace_tree_ w111(.clk(clk),.rst_n(rst_n),.a({x_0[111],x_1[111],x_2[111],x_3[111],x_4[111],x_5[111],x_6[111],x_7[111],x_8[111],x_9[111],x_10[111],x_11[111],x_12[111],x_13[111],x_14[111],x_15[111],x_16[111],x_17[111],x_18[111],x_19[111],x_20[111],x_21[111],x_22[111],x_23[111],x_24[111],x_25[111],x_26[111],x_27[111],x_28[111],x_29[111],x_30[111],x_31[111],x_32[111]}),.c_in(c_in_111),.c_out(c_in_112),.s(s_111),.c(c_111));
wire  c_112;
wire  s_112;
wallace_tree_ w112(.clk(clk),.rst_n(rst_n),.a({x_0[112],x_1[112],x_2[112],x_3[112],x_4[112],x_5[112],x_6[112],x_7[112],x_8[112],x_9[112],x_10[112],x_11[112],x_12[112],x_13[112],x_14[112],x_15[112],x_16[112],x_17[112],x_18[112],x_19[112],x_20[112],x_21[112],x_22[112],x_23[112],x_24[112],x_25[112],x_26[112],x_27[112],x_28[112],x_29[112],x_30[112],x_31[112],x_32[112]}),.c_in(c_in_112),.c_out(c_in_113),.s(s_112),.c(c_112));
wire  c_113;
wire  s_113;
wallace_tree_ w113(.clk(clk),.rst_n(rst_n),.a({x_0[113],x_1[113],x_2[113],x_3[113],x_4[113],x_5[113],x_6[113],x_7[113],x_8[113],x_9[113],x_10[113],x_11[113],x_12[113],x_13[113],x_14[113],x_15[113],x_16[113],x_17[113],x_18[113],x_19[113],x_20[113],x_21[113],x_22[113],x_23[113],x_24[113],x_25[113],x_26[113],x_27[113],x_28[113],x_29[113],x_30[113],x_31[113],x_32[113]}),.c_in(c_in_113),.c_out(c_in_114),.s(s_113),.c(c_113));
wire  c_114;
wire  s_114;
wallace_tree_ w114(.clk(clk),.rst_n(rst_n),.a({x_0[114],x_1[114],x_2[114],x_3[114],x_4[114],x_5[114],x_6[114],x_7[114],x_8[114],x_9[114],x_10[114],x_11[114],x_12[114],x_13[114],x_14[114],x_15[114],x_16[114],x_17[114],x_18[114],x_19[114],x_20[114],x_21[114],x_22[114],x_23[114],x_24[114],x_25[114],x_26[114],x_27[114],x_28[114],x_29[114],x_30[114],x_31[114],x_32[114]}),.c_in(c_in_114),.c_out(c_in_115),.s(s_114),.c(c_114));
wire  c_115;
wire  s_115;
wallace_tree_ w115(.clk(clk),.rst_n(rst_n),.a({x_0[115],x_1[115],x_2[115],x_3[115],x_4[115],x_5[115],x_6[115],x_7[115],x_8[115],x_9[115],x_10[115],x_11[115],x_12[115],x_13[115],x_14[115],x_15[115],x_16[115],x_17[115],x_18[115],x_19[115],x_20[115],x_21[115],x_22[115],x_23[115],x_24[115],x_25[115],x_26[115],x_27[115],x_28[115],x_29[115],x_30[115],x_31[115],x_32[115]}),.c_in(c_in_115),.c_out(c_in_116),.s(s_115),.c(c_115));
wire  c_116;
wire  s_116;
wallace_tree_ w116(.clk(clk),.rst_n(rst_n),.a({x_0[116],x_1[116],x_2[116],x_3[116],x_4[116],x_5[116],x_6[116],x_7[116],x_8[116],x_9[116],x_10[116],x_11[116],x_12[116],x_13[116],x_14[116],x_15[116],x_16[116],x_17[116],x_18[116],x_19[116],x_20[116],x_21[116],x_22[116],x_23[116],x_24[116],x_25[116],x_26[116],x_27[116],x_28[116],x_29[116],x_30[116],x_31[116],x_32[116]}),.c_in(c_in_116),.c_out(c_in_117),.s(s_116),.c(c_116));
wire  c_117;
wire  s_117;
wallace_tree_ w117(.clk(clk),.rst_n(rst_n),.a({x_0[117],x_1[117],x_2[117],x_3[117],x_4[117],x_5[117],x_6[117],x_7[117],x_8[117],x_9[117],x_10[117],x_11[117],x_12[117],x_13[117],x_14[117],x_15[117],x_16[117],x_17[117],x_18[117],x_19[117],x_20[117],x_21[117],x_22[117],x_23[117],x_24[117],x_25[117],x_26[117],x_27[117],x_28[117],x_29[117],x_30[117],x_31[117],x_32[117]}),.c_in(c_in_117),.c_out(c_in_118),.s(s_117),.c(c_117));
wire  c_118;
wire  s_118;
wallace_tree_ w118(.clk(clk),.rst_n(rst_n),.a({x_0[118],x_1[118],x_2[118],x_3[118],x_4[118],x_5[118],x_6[118],x_7[118],x_8[118],x_9[118],x_10[118],x_11[118],x_12[118],x_13[118],x_14[118],x_15[118],x_16[118],x_17[118],x_18[118],x_19[118],x_20[118],x_21[118],x_22[118],x_23[118],x_24[118],x_25[118],x_26[118],x_27[118],x_28[118],x_29[118],x_30[118],x_31[118],x_32[118]}),.c_in(c_in_118),.c_out(c_in_119),.s(s_118),.c(c_118));
wire  c_119;
wire  s_119;
wallace_tree_ w119(.clk(clk),.rst_n(rst_n),.a({x_0[119],x_1[119],x_2[119],x_3[119],x_4[119],x_5[119],x_6[119],x_7[119],x_8[119],x_9[119],x_10[119],x_11[119],x_12[119],x_13[119],x_14[119],x_15[119],x_16[119],x_17[119],x_18[119],x_19[119],x_20[119],x_21[119],x_22[119],x_23[119],x_24[119],x_25[119],x_26[119],x_27[119],x_28[119],x_29[119],x_30[119],x_31[119],x_32[119]}),.c_in(c_in_119),.c_out(c_in_120),.s(s_119),.c(c_119));
wire  c_120;
wire  s_120;
wallace_tree_ w120(.clk(clk),.rst_n(rst_n),.a({x_0[120],x_1[120],x_2[120],x_3[120],x_4[120],x_5[120],x_6[120],x_7[120],x_8[120],x_9[120],x_10[120],x_11[120],x_12[120],x_13[120],x_14[120],x_15[120],x_16[120],x_17[120],x_18[120],x_19[120],x_20[120],x_21[120],x_22[120],x_23[120],x_24[120],x_25[120],x_26[120],x_27[120],x_28[120],x_29[120],x_30[120],x_31[120],x_32[120]}),.c_in(c_in_120),.c_out(c_in_121),.s(s_120),.c(c_120));
wire  c_121;
wire  s_121;
wallace_tree_ w121(.clk(clk),.rst_n(rst_n),.a({x_0[121],x_1[121],x_2[121],x_3[121],x_4[121],x_5[121],x_6[121],x_7[121],x_8[121],x_9[121],x_10[121],x_11[121],x_12[121],x_13[121],x_14[121],x_15[121],x_16[121],x_17[121],x_18[121],x_19[121],x_20[121],x_21[121],x_22[121],x_23[121],x_24[121],x_25[121],x_26[121],x_27[121],x_28[121],x_29[121],x_30[121],x_31[121],x_32[121]}),.c_in(c_in_121),.c_out(c_in_122),.s(s_121),.c(c_121));
wire  c_122;
wire  s_122;
wallace_tree_ w122(.clk(clk),.rst_n(rst_n),.a({x_0[122],x_1[122],x_2[122],x_3[122],x_4[122],x_5[122],x_6[122],x_7[122],x_8[122],x_9[122],x_10[122],x_11[122],x_12[122],x_13[122],x_14[122],x_15[122],x_16[122],x_17[122],x_18[122],x_19[122],x_20[122],x_21[122],x_22[122],x_23[122],x_24[122],x_25[122],x_26[122],x_27[122],x_28[122],x_29[122],x_30[122],x_31[122],x_32[122]}),.c_in(c_in_122),.c_out(c_in_123),.s(s_122),.c(c_122));
wire  c_123;
wire  s_123;
wallace_tree_ w123(.clk(clk),.rst_n(rst_n),.a({x_0[123],x_1[123],x_2[123],x_3[123],x_4[123],x_5[123],x_6[123],x_7[123],x_8[123],x_9[123],x_10[123],x_11[123],x_12[123],x_13[123],x_14[123],x_15[123],x_16[123],x_17[123],x_18[123],x_19[123],x_20[123],x_21[123],x_22[123],x_23[123],x_24[123],x_25[123],x_26[123],x_27[123],x_28[123],x_29[123],x_30[123],x_31[123],x_32[123]}),.c_in(c_in_123),.c_out(c_in_124),.s(s_123),.c(c_123));
wire  c_124;
wire  s_124;
wallace_tree_ w124(.clk(clk),.rst_n(rst_n),.a({x_0[124],x_1[124],x_2[124],x_3[124],x_4[124],x_5[124],x_6[124],x_7[124],x_8[124],x_9[124],x_10[124],x_11[124],x_12[124],x_13[124],x_14[124],x_15[124],x_16[124],x_17[124],x_18[124],x_19[124],x_20[124],x_21[124],x_22[124],x_23[124],x_24[124],x_25[124],x_26[124],x_27[124],x_28[124],x_29[124],x_30[124],x_31[124],x_32[124]}),.c_in(c_in_124),.c_out(c_in_125),.s(s_124),.c(c_124));
wire  c_125;
wire  s_125;
wallace_tree_ w125(.clk(clk),.rst_n(rst_n),.a({x_0[125],x_1[125],x_2[125],x_3[125],x_4[125],x_5[125],x_6[125],x_7[125],x_8[125],x_9[125],x_10[125],x_11[125],x_12[125],x_13[125],x_14[125],x_15[125],x_16[125],x_17[125],x_18[125],x_19[125],x_20[125],x_21[125],x_22[125],x_23[125],x_24[125],x_25[125],x_26[125],x_27[125],x_28[125],x_29[125],x_30[125],x_31[125],x_32[125]}),.c_in(c_in_125),.c_out(c_in_126),.s(s_125),.c(c_125));
wire  c_126;
wire  s_126;
wallace_tree_ w126(.clk(clk),.rst_n(rst_n),.a({x_0[126],x_1[126],x_2[126],x_3[126],x_4[126],x_5[126],x_6[126],x_7[126],x_8[126],x_9[126],x_10[126],x_11[126],x_12[126],x_13[126],x_14[126],x_15[126],x_16[126],x_17[126],x_18[126],x_19[126],x_20[126],x_21[126],x_22[126],x_23[126],x_24[126],x_25[126],x_26[126],x_27[126],x_28[126],x_29[126],x_30[126],x_31[126],x_32[126]}),.c_in(c_in_126),.c_out(c_in_127),.s(s_126),.c(c_126));
wire  c_127;
wire  s_127;
wallace_tree_ w127(.clk(clk),.rst_n(rst_n),.a({x_0[127],x_1[127],x_2[127],x_3[127],x_4[127],x_5[127],x_6[127],x_7[127],x_8[127],x_9[127],x_10[127],x_11[127],x_12[127],x_13[127],x_14[127],x_15[127],x_16[127],x_17[127],x_18[127],x_19[127],x_20[127],x_21[127],x_22[127],x_23[127],x_24[127],x_25[127],x_26[127],x_27[127],x_28[127],x_29[127],x_30[127],x_31[127],x_32[127]}),.c_in(c_in_127),.c_out(c_in_128),.s(s_127),.c(c_127));
wire  c_128;
wire  s_128;
wallace_tree_ w128(.clk(clk),.rst_n(rst_n),.a({x_0[128],x_1[128],x_2[128],x_3[128],x_4[128],x_5[128],x_6[128],x_7[128],x_8[128],x_9[128],x_10[128],x_11[128],x_12[128],x_13[128],x_14[128],x_15[128],x_16[128],x_17[128],x_18[128],x_19[128],x_20[128],x_21[128],x_22[128],x_23[128],x_24[128],x_25[128],x_26[128],x_27[128],x_28[128],x_29[128],x_30[128],x_31[128],x_32[128]}),.c_in(c_in_128),.c_out(c_in_129),.s(s_128),.c(c_128));
wire  c_129;
wire  s_129;
wallace_tree_ w129(.clk(clk),.rst_n(rst_n),.a({x_0[129],x_1[129],x_2[129],x_3[129],x_4[129],x_5[129],x_6[129],x_7[129],x_8[129],x_9[129],x_10[129],x_11[129],x_12[129],x_13[129],x_14[129],x_15[129],x_16[129],x_17[129],x_18[129],x_19[129],x_20[129],x_21[129],x_22[129],x_23[129],x_24[129],x_25[129],x_26[129],x_27[129],x_28[129],x_29[129],x_30[129],x_31[129],x_32[129]}),.c_in(c_in_129),.c_out(c_in_130),.s(s_129),.c(c_129));
wire  c_130;
wire  s_130;
wallace_tree_ w130(.clk(clk),.rst_n(rst_n),.a({x_0[130],x_1[130],x_2[130],x_3[130],x_4[130],x_5[130],x_6[130],x_7[130],x_8[130],x_9[130],x_10[130],x_11[130],x_12[130],x_13[130],x_14[130],x_15[130],x_16[130],x_17[130],x_18[130],x_19[130],x_20[130],x_21[130],x_22[130],x_23[130],x_24[130],x_25[130],x_26[130],x_27[130],x_28[130],x_29[130],x_30[130],x_31[130],x_32[130]}),.c_in(c_in_130),.c_out(c_in_131),.s(s_130),.c(c_130));
wire  c_131;
wire  s_131;
wallace_tree_ w131(.clk(clk),.rst_n(rst_n),.a({x_0[131],x_1[131],x_2[131],x_3[131],x_4[131],x_5[131],x_6[131],x_7[131],x_8[131],x_9[131],x_10[131],x_11[131],x_12[131],x_13[131],x_14[131],x_15[131],x_16[131],x_17[131],x_18[131],x_19[131],x_20[131],x_21[131],x_22[131],x_23[131],x_24[131],x_25[131],x_26[131],x_27[131],x_28[131],x_29[131],x_30[131],x_31[131],x_32[131]}),.c_in(c_in_131),.c_out(),.s(s_131),.c(c_131));
assign s = {s_131,s_130,s_129,s_128,s_127,s_126,s_125,s_124,s_123,s_122,s_121,s_120,s_119,s_118,s_117,s_116,s_115,s_114,s_113,s_112,s_111,s_110,s_109,s_108,s_107,s_106,s_105,s_104,s_103,s_102,s_101,s_100,s_99,s_98,s_97,s_96,s_95,s_94,s_93,s_92,s_91,s_90,s_89,s_88,s_87,s_86,s_85,s_84,s_83,s_82,s_81,s_80,s_79,s_78,s_77,s_76,s_75,s_74,s_73,s_72,s_71,s_70,s_69,s_68,s_67,s_66,s_65,s_64,s_63,s_62,s_61,s_60,s_59,s_58,s_57,s_56,s_55,s_54,s_53,s_52,s_51,s_50,s_49,s_48,s_47,s_46,s_45,s_44,s_43,s_42,s_41,s_40,s_39,s_38,s_37,s_36,s_35,s_34,s_33,s_32,s_31,s_30,s_29,s_28,s_27,s_26,s_25,s_24,s_23,s_22,s_21,s_20,s_19,s_18,s_17,s_16,s_15,s_14,s_13,s_12,s_11,s_10,s_9,s_8,s_7,s_6,s_5,s_4,s_3,s_2,s_1,s_0 };
assign c = {c_131,c_130,c_129,c_128,c_127,c_126,c_125,c_124,c_123,c_122,c_121,c_120,c_119,c_118,c_117,c_116,c_115,c_114,c_113,c_112,c_111,c_110,c_109,c_108,c_107,c_106,c_105,c_104,c_103,c_102,c_101,c_100,c_99,c_98,c_97,c_96,c_95,c_94,c_93,c_92,c_91,c_90,c_89,c_88,c_87,c_86,c_85,c_84,c_83,c_82,c_81,c_80,c_79,c_78,c_77,c_76,c_75,c_74,c_73,c_72,c_71,c_70,c_69,c_68,c_67,c_66,c_65,c_64,c_63,c_62,c_61,c_60,c_59,c_58,c_57,c_56,c_55,c_54,c_53,c_52,c_51,c_50,c_49,c_48,c_47,c_46,c_45,c_44,c_43,c_42,c_41,c_40,c_39,c_38,c_37,c_36,c_35,c_34,c_33,c_32,c_31,c_30,c_29,c_28,c_27,c_26,c_25,c_24,c_23,c_22,c_21,c_20,c_19,c_18,c_17,c_16,c_15,c_14,c_13,c_12,c_11,c_10,c_9,c_8,c_7,c_6,c_5,c_4,c_3,c_2,c_1,c_0 };
endmodule