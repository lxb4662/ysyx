module ysyx_22050518_add (
 input [63:0]    in1, 
 input [63:0]    in2,
 input              c_in,
 output [63:0]    out 
);
 wire [63:0]    a;
 wire [63:0]    b;
 wire [63:0]    g;
 wire [63:0]    p;
  wire [63:0]    s;
assign c_0 = c_in;
assign a = in1;
assign b = in2;
wire c_0; 
wire c_1; 
wire c_2; 
wire c_3; 
wire c_4; 
wire c_5; 
wire c_6; 
wire c_7; 
wire c_8; 
wire c_9; 
wire c_10; 
wire c_11; 
wire c_12; 
wire c_13; 
wire c_14; 
wire c_15; 
wire c_16; 
wire c_17; 
wire c_18; 
wire c_19; 
wire c_20; 
wire c_21; 
wire c_22; 
wire c_23; 
wire c_24; 
wire c_25; 
wire c_26; 
wire c_27; 
wire c_28; 
wire c_29; 
wire c_30; 
wire c_31; 
wire c_32; 
wire c_33; 
wire c_34; 
wire c_35; 
wire c_36; 
wire c_37; 
wire c_38; 
wire c_39; 
wire c_40; 
wire c_41; 
wire c_42; 
wire c_43; 
wire c_44; 
wire c_45; 
wire c_46; 
wire c_47; 
wire c_48; 
wire c_49; 
wire c_50; 
wire c_51; 
wire c_52; 
wire c_53; 
wire c_54; 
wire c_55; 
wire c_56; 
wire c_57; 
wire c_58; 
wire c_59; 
wire c_60; 
wire c_61; 
wire c_62; 
wire c_63; 
full_adder_1bit full_adder_0(.a(a[0]),.b(b[0]),.c_in(c_0),.c_out(),.s(s[0]));
full_adder_1bit full_adder_1(.a(a[1]),.b(b[1]),.c_in(c_1),.c_out(),.s(s[1]));
full_adder_1bit full_adder_2(.a(a[2]),.b(b[2]),.c_in(c_2),.c_out(),.s(s[2]));
full_adder_1bit full_adder_3(.a(a[3]),.b(b[3]),.c_in(c_3),.c_out(),.s(s[3]));
full_adder_1bit full_adder_4(.a(a[4]),.b(b[4]),.c_in(c_4),.c_out(),.s(s[4]));
full_adder_1bit full_adder_5(.a(a[5]),.b(b[5]),.c_in(c_5),.c_out(),.s(s[5]));
full_adder_1bit full_adder_6(.a(a[6]),.b(b[6]),.c_in(c_6),.c_out(),.s(s[6]));
full_adder_1bit full_adder_7(.a(a[7]),.b(b[7]),.c_in(c_7),.c_out(),.s(s[7]));
full_adder_1bit full_adder_8(.a(a[8]),.b(b[8]),.c_in(c_8),.c_out(),.s(s[8]));
full_adder_1bit full_adder_9(.a(a[9]),.b(b[9]),.c_in(c_9),.c_out(),.s(s[9]));
full_adder_1bit full_adder_10(.a(a[10]),.b(b[10]),.c_in(c_10),.c_out(),.s(s[10]));
full_adder_1bit full_adder_11(.a(a[11]),.b(b[11]),.c_in(c_11),.c_out(),.s(s[11]));
full_adder_1bit full_adder_12(.a(a[12]),.b(b[12]),.c_in(c_12),.c_out(),.s(s[12]));
full_adder_1bit full_adder_13(.a(a[13]),.b(b[13]),.c_in(c_13),.c_out(),.s(s[13]));
full_adder_1bit full_adder_14(.a(a[14]),.b(b[14]),.c_in(c_14),.c_out(),.s(s[14]));
full_adder_1bit full_adder_15(.a(a[15]),.b(b[15]),.c_in(c_15),.c_out(),.s(s[15]));
full_adder_1bit full_adder_16(.a(a[16]),.b(b[16]),.c_in(c_16),.c_out(),.s(s[16]));
full_adder_1bit full_adder_17(.a(a[17]),.b(b[17]),.c_in(c_17),.c_out(),.s(s[17]));
full_adder_1bit full_adder_18(.a(a[18]),.b(b[18]),.c_in(c_18),.c_out(),.s(s[18]));
full_adder_1bit full_adder_19(.a(a[19]),.b(b[19]),.c_in(c_19),.c_out(),.s(s[19]));
full_adder_1bit full_adder_20(.a(a[20]),.b(b[20]),.c_in(c_20),.c_out(),.s(s[20]));
full_adder_1bit full_adder_21(.a(a[21]),.b(b[21]),.c_in(c_21),.c_out(),.s(s[21]));
full_adder_1bit full_adder_22(.a(a[22]),.b(b[22]),.c_in(c_22),.c_out(),.s(s[22]));
full_adder_1bit full_adder_23(.a(a[23]),.b(b[23]),.c_in(c_23),.c_out(),.s(s[23]));
full_adder_1bit full_adder_24(.a(a[24]),.b(b[24]),.c_in(c_24),.c_out(),.s(s[24]));
full_adder_1bit full_adder_25(.a(a[25]),.b(b[25]),.c_in(c_25),.c_out(),.s(s[25]));
full_adder_1bit full_adder_26(.a(a[26]),.b(b[26]),.c_in(c_26),.c_out(),.s(s[26]));
full_adder_1bit full_adder_27(.a(a[27]),.b(b[27]),.c_in(c_27),.c_out(),.s(s[27]));
full_adder_1bit full_adder_28(.a(a[28]),.b(b[28]),.c_in(c_28),.c_out(),.s(s[28]));
full_adder_1bit full_adder_29(.a(a[29]),.b(b[29]),.c_in(c_29),.c_out(),.s(s[29]));
full_adder_1bit full_adder_30(.a(a[30]),.b(b[30]),.c_in(c_30),.c_out(),.s(s[30]));
full_adder_1bit full_adder_31(.a(a[31]),.b(b[31]),.c_in(c_31),.c_out(),.s(s[31]));
full_adder_1bit full_adder_32(.a(a[32]),.b(b[32]),.c_in(c_32),.c_out(),.s(s[32]));
full_adder_1bit full_adder_33(.a(a[33]),.b(b[33]),.c_in(c_33),.c_out(),.s(s[33]));
full_adder_1bit full_adder_34(.a(a[34]),.b(b[34]),.c_in(c_34),.c_out(),.s(s[34]));
full_adder_1bit full_adder_35(.a(a[35]),.b(b[35]),.c_in(c_35),.c_out(),.s(s[35]));
full_adder_1bit full_adder_36(.a(a[36]),.b(b[36]),.c_in(c_36),.c_out(),.s(s[36]));
full_adder_1bit full_adder_37(.a(a[37]),.b(b[37]),.c_in(c_37),.c_out(),.s(s[37]));
full_adder_1bit full_adder_38(.a(a[38]),.b(b[38]),.c_in(c_38),.c_out(),.s(s[38]));
full_adder_1bit full_adder_39(.a(a[39]),.b(b[39]),.c_in(c_39),.c_out(),.s(s[39]));
full_adder_1bit full_adder_40(.a(a[40]),.b(b[40]),.c_in(c_40),.c_out(),.s(s[40]));
full_adder_1bit full_adder_41(.a(a[41]),.b(b[41]),.c_in(c_41),.c_out(),.s(s[41]));
full_adder_1bit full_adder_42(.a(a[42]),.b(b[42]),.c_in(c_42),.c_out(),.s(s[42]));
full_adder_1bit full_adder_43(.a(a[43]),.b(b[43]),.c_in(c_43),.c_out(),.s(s[43]));
full_adder_1bit full_adder_44(.a(a[44]),.b(b[44]),.c_in(c_44),.c_out(),.s(s[44]));
full_adder_1bit full_adder_45(.a(a[45]),.b(b[45]),.c_in(c_45),.c_out(),.s(s[45]));
full_adder_1bit full_adder_46(.a(a[46]),.b(b[46]),.c_in(c_46),.c_out(),.s(s[46]));
full_adder_1bit full_adder_47(.a(a[47]),.b(b[47]),.c_in(c_47),.c_out(),.s(s[47]));
full_adder_1bit full_adder_48(.a(a[48]),.b(b[48]),.c_in(c_48),.c_out(),.s(s[48]));
full_adder_1bit full_adder_49(.a(a[49]),.b(b[49]),.c_in(c_49),.c_out(),.s(s[49]));
full_adder_1bit full_adder_50(.a(a[50]),.b(b[50]),.c_in(c_50),.c_out(),.s(s[50]));
full_adder_1bit full_adder_51(.a(a[51]),.b(b[51]),.c_in(c_51),.c_out(),.s(s[51]));
full_adder_1bit full_adder_52(.a(a[52]),.b(b[52]),.c_in(c_52),.c_out(),.s(s[52]));
full_adder_1bit full_adder_53(.a(a[53]),.b(b[53]),.c_in(c_53),.c_out(),.s(s[53]));
full_adder_1bit full_adder_54(.a(a[54]),.b(b[54]),.c_in(c_54),.c_out(),.s(s[54]));
full_adder_1bit full_adder_55(.a(a[55]),.b(b[55]),.c_in(c_55),.c_out(),.s(s[55]));
full_adder_1bit full_adder_56(.a(a[56]),.b(b[56]),.c_in(c_56),.c_out(),.s(s[56]));
full_adder_1bit full_adder_57(.a(a[57]),.b(b[57]),.c_in(c_57),.c_out(),.s(s[57]));
full_adder_1bit full_adder_58(.a(a[58]),.b(b[58]),.c_in(c_58),.c_out(),.s(s[58]));
full_adder_1bit full_adder_59(.a(a[59]),.b(b[59]),.c_in(c_59),.c_out(),.s(s[59]));
full_adder_1bit full_adder_60(.a(a[60]),.b(b[60]),.c_in(c_60),.c_out(),.s(s[60]));
full_adder_1bit full_adder_61(.a(a[61]),.b(b[61]),.c_in(c_61),.c_out(),.s(s[61]));
full_adder_1bit full_adder_62(.a(a[62]),.b(b[62]),.c_in(c_62),.c_out(),.s(s[62]));
full_adder_1bit full_adder_63(.a(a[63]),.b(b[63]),.c_in(c_63),.c_out(),.s(s[63]));
assign g[0]    = a[0]&b[0];
assign p[0]    = a[0]|b[0];
assign c_1    = g[0]|p[0]&c_0;
assign g[1]    = a[1]&b[1];
assign p[1]    = a[1]|b[1];
assign c_2    = g[1]|p[1]&c_1;
assign g[2]    = a[2]&b[2];
assign p[2]    = a[2]|b[2];
assign c_3    = g[2]|p[2]&c_2;
assign g[3]    = a[3]&b[3];
assign p[3]    = a[3]|b[3];
assign c_4    = g[3]|p[3]&c_3;
assign g[4]    = a[4]&b[4];
assign p[4]    = a[4]|b[4];
assign c_5    = g[4]|p[4]&c_4;
assign g[5]    = a[5]&b[5];
assign p[5]    = a[5]|b[5];
assign c_6    = g[5]|p[5]&c_5;
assign g[6]    = a[6]&b[6];
assign p[6]    = a[6]|b[6];
assign c_7    = g[6]|p[6]&c_6;
assign g[7]    = a[7]&b[7];
assign p[7]    = a[7]|b[7];
assign c_8    = g[7]|p[7]&c_7;
assign g[8]    = a[8]&b[8];
assign p[8]    = a[8]|b[8];
assign c_9    = g[8]|p[8]&c_8;
assign g[9]    = a[9]&b[9];
assign p[9]    = a[9]|b[9];
assign c_10    = g[9]|p[9]&c_9;
assign g[10]    = a[10]&b[10];
assign p[10]    = a[10]|b[10];
assign c_11    = g[10]|p[10]&c_10;
assign g[11]    = a[11]&b[11];
assign p[11]    = a[11]|b[11];
assign c_12    = g[11]|p[11]&c_11;
assign g[12]    = a[12]&b[12];
assign p[12]    = a[12]|b[12];
assign c_13    = g[12]|p[12]&c_12;
assign g[13]    = a[13]&b[13];
assign p[13]    = a[13]|b[13];
assign c_14    = g[13]|p[13]&c_13;
assign g[14]    = a[14]&b[14];
assign p[14]    = a[14]|b[14];
assign c_15    = g[14]|p[14]&c_14;
assign g[15]    = a[15]&b[15];
assign p[15]    = a[15]|b[15];
assign c_16    = g[15]|p[15]&c_15;
assign g[16]    = a[16]&b[16];
assign p[16]    = a[16]|b[16];
assign c_17    = g[16]|p[16]&c_16;
assign g[17]    = a[17]&b[17];
assign p[17]    = a[17]|b[17];
assign c_18    = g[17]|p[17]&c_17;
assign g[18]    = a[18]&b[18];
assign p[18]    = a[18]|b[18];
assign c_19    = g[18]|p[18]&c_18;
assign g[19]    = a[19]&b[19];
assign p[19]    = a[19]|b[19];
assign c_20    = g[19]|p[19]&c_19;
assign g[20]    = a[20]&b[20];
assign p[20]    = a[20]|b[20];
assign c_21    = g[20]|p[20]&c_20;
assign g[21]    = a[21]&b[21];
assign p[21]    = a[21]|b[21];
assign c_22    = g[21]|p[21]&c_21;
assign g[22]    = a[22]&b[22];
assign p[22]    = a[22]|b[22];
assign c_23    = g[22]|p[22]&c_22;
assign g[23]    = a[23]&b[23];
assign p[23]    = a[23]|b[23];
assign c_24    = g[23]|p[23]&c_23;
assign g[24]    = a[24]&b[24];
assign p[24]    = a[24]|b[24];
assign c_25    = g[24]|p[24]&c_24;
assign g[25]    = a[25]&b[25];
assign p[25]    = a[25]|b[25];
assign c_26    = g[25]|p[25]&c_25;
assign g[26]    = a[26]&b[26];
assign p[26]    = a[26]|b[26];
assign c_27    = g[26]|p[26]&c_26;
assign g[27]    = a[27]&b[27];
assign p[27]    = a[27]|b[27];
assign c_28    = g[27]|p[27]&c_27;
assign g[28]    = a[28]&b[28];
assign p[28]    = a[28]|b[28];
assign c_29    = g[28]|p[28]&c_28;
assign g[29]    = a[29]&b[29];
assign p[29]    = a[29]|b[29];
assign c_30    = g[29]|p[29]&c_29;
assign g[30]    = a[30]&b[30];
assign p[30]    = a[30]|b[30];
assign c_31    = g[30]|p[30]&c_30;
assign g[31]    = a[31]&b[31];
assign p[31]    = a[31]|b[31];
assign c_32    = g[31]|p[31]&c_31;
assign g[32]    = a[32]&b[32];
assign p[32]    = a[32]|b[32];
assign c_33    = g[32]|p[32]&c_32;
assign g[33]    = a[33]&b[33];
assign p[33]    = a[33]|b[33];
assign c_34    = g[33]|p[33]&c_33;
assign g[34]    = a[34]&b[34];
assign p[34]    = a[34]|b[34];
assign c_35    = g[34]|p[34]&c_34;
assign g[35]    = a[35]&b[35];
assign p[35]    = a[35]|b[35];
assign c_36    = g[35]|p[35]&c_35;
assign g[36]    = a[36]&b[36];
assign p[36]    = a[36]|b[36];
assign c_37    = g[36]|p[36]&c_36;
assign g[37]    = a[37]&b[37];
assign p[37]    = a[37]|b[37];
assign c_38    = g[37]|p[37]&c_37;
assign g[38]    = a[38]&b[38];
assign p[38]    = a[38]|b[38];
assign c_39    = g[38]|p[38]&c_38;
assign g[39]    = a[39]&b[39];
assign p[39]    = a[39]|b[39];
assign c_40    = g[39]|p[39]&c_39;
assign g[40]    = a[40]&b[40];
assign p[40]    = a[40]|b[40];
assign c_41    = g[40]|p[40]&c_40;
assign g[41]    = a[41]&b[41];
assign p[41]    = a[41]|b[41];
assign c_42    = g[41]|p[41]&c_41;
assign g[42]    = a[42]&b[42];
assign p[42]    = a[42]|b[42];
assign c_43    = g[42]|p[42]&c_42;
assign g[43]    = a[43]&b[43];
assign p[43]    = a[43]|b[43];
assign c_44    = g[43]|p[43]&c_43;
assign g[44]    = a[44]&b[44];
assign p[44]    = a[44]|b[44];
assign c_45    = g[44]|p[44]&c_44;
assign g[45]    = a[45]&b[45];
assign p[45]    = a[45]|b[45];
assign c_46    = g[45]|p[45]&c_45;
assign g[46]    = a[46]&b[46];
assign p[46]    = a[46]|b[46];
assign c_47    = g[46]|p[46]&c_46;
assign g[47]    = a[47]&b[47];
assign p[47]    = a[47]|b[47];
assign c_48    = g[47]|p[47]&c_47;
assign g[48]    = a[48]&b[48];
assign p[48]    = a[48]|b[48];
assign c_49    = g[48]|p[48]&c_48;
assign g[49]    = a[49]&b[49];
assign p[49]    = a[49]|b[49];
assign c_50    = g[49]|p[49]&c_49;
assign g[50]    = a[50]&b[50];
assign p[50]    = a[50]|b[50];
assign c_51    = g[50]|p[50]&c_50;
assign g[51]    = a[51]&b[51];
assign p[51]    = a[51]|b[51];
assign c_52    = g[51]|p[51]&c_51;
assign g[52]    = a[52]&b[52];
assign p[52]    = a[52]|b[52];
assign c_53    = g[52]|p[52]&c_52;
assign g[53]    = a[53]&b[53];
assign p[53]    = a[53]|b[53];
assign c_54    = g[53]|p[53]&c_53;
assign g[54]    = a[54]&b[54];
assign p[54]    = a[54]|b[54];
assign c_55    = g[54]|p[54]&c_54;
assign g[55]    = a[55]&b[55];
assign p[55]    = a[55]|b[55];
assign c_56    = g[55]|p[55]&c_55;
assign g[56]    = a[56]&b[56];
assign p[56]    = a[56]|b[56];
assign c_57    = g[56]|p[56]&c_56;
assign g[57]    = a[57]&b[57];
assign p[57]    = a[57]|b[57];
assign c_58    = g[57]|p[57]&c_57;
assign g[58]    = a[58]&b[58];
assign p[58]    = a[58]|b[58];
assign c_59    = g[58]|p[58]&c_58;
assign g[59]    = a[59]&b[59];
assign p[59]    = a[59]|b[59];
assign c_60    = g[59]|p[59]&c_59;
assign g[60]    = a[60]&b[60];
assign p[60]    = a[60]|b[60];
assign c_61    = g[60]|p[60]&c_60;
assign g[61]    = a[61]&b[61];
assign p[61]    = a[61]|b[61];
assign c_62    = g[61]|p[61]&c_61;
assign g[62]    = a[62]&b[62];
assign p[62]    = a[62]|b[62];
assign c_63    = g[62]|p[62]&c_62;
assign g[63]    = a[63]&b[63];
assign p[63]    = a[63]|b[63];
//assign c_64    = g[63]|p[63]&c_63;
assign out = s;
endmodule 

